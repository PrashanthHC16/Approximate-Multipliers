-- Owner : Prashanth H C,( prashanth.c@iiitb.ac.in )
-- File part of SOMALib Activation functions library
-- All circuits : https://github.com/PrashanthHC16/Activation-Functions-Library
-- The file is distributed under MIT License.


LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY tanh_Config2_Approx_10_4bit_B_cir2 IS
PORT( Inp                               :   IN    std_logic_vector(3 downto 0);
      Out1                             :   OUT   std_logic_vector(3 downto 0)
      );
END tanh_Config2_Approx_10_4bit_B_cir2;


ARCHITECTURE rtl OF tanh_Config2_Approx_10_4bit_B_cir2 IS

-- Signals
SIGNAL XOR0_out1                        : std_logic;
SIGNAL XOR4_out1                        : std_logic;
SIGNAL NOR2_out1                        : std_logic;
SIGNAL NAND1_out1                       : std_logic;
SIGNAL AND3_out1                        : std_logic;
SIGNAL NOR5_out1                        : std_logic;

BEGIN
XOR0_out1 <= Inp(0) XOR Inp(2);

XOR4_out1 <= Inp(2) XOR XOR0_out1;

NOR2_out1 <=  NOT (XOR0_out1 OR Inp(1));

NAND1_out1 <=  NOT (Inp(2) AND Inp(3));

AND3_out1 <= Inp(0) AND NAND1_out1;

NOR5_out1 <=  NOT (NOR2_out1 OR AND3_out1);

Out1(0) <= XOR4_out1;

Out1(1) <= XOR4_out1;

Out1(2) <= NOR5_out1;

Out1(3) <= NOR5_out1;

END rtl;
