///////////////////////////////////////////////////////////////////////////////////////////////////
// Owned by : Prashanth H C, Prashanth.C@iiitb.ac.in / prashanth.c@iiitb.org
// File distributed under MIT License.
// 2021 September
//
// Complete implementation : https://github.com/PrashanthHC16/Approximate-Multipliers
//
// Part of paper "Performance and Error Analysis of Approximate Multipliers of Different Configurations and Fast Adders"
// Authors : Prashanth H C, Soujanya S R, Bindu G Gowda, Madhav Rao
//
///////////////////////////////////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps


module dadda_processing_block_16(  // Owner : Soujanya S R, soujanya.sr@iiitb.ac.in 
        input    pp [15:0][15:0],
        output [31:0] to_FA [1:0]      
    );
    //requires 195 FA;
    //requies 15 HA
    
    //#of full adder sum & carry to be captured
    //195 - 27 = 168 reg required for each as last set o/p will be directly connected to the o/p
    reg fs[167:0];
    reg fc[167:0];
    
    //15-1 = 14 reg required
    reg hs[13:0];
    reg hc[13:0];
    
  /////////////////////////////// RS1 16 -> 13 /////////////////////////////////
  // Adders: FA = 8; HA = 4
  
  fa fa0  (.A(pp[00][14]), .B(pp[01][13]), .Ci(pp[02][12]), .S(fs[0]), .Co(fc[0]));
  fa fa1  (.A(pp[00][15]), .B(pp[01][14]), .Ci(pp[02][13]), .S(fs[1]), .Co(fc[1]));
  fa fa2  (.A(pp[03][12]), .B(pp[04][11]), .Ci(pp[05][10]), .S(fs[2]), .Co(fc[2]));
  fa fa3  (.A(pp[01][15]), .B(pp[02][14]), .Ci(pp[03][13]), .S(fs[3]), .Co(fc[3]));
  fa fa4  (.A(pp[04][12]), .B(pp[05][11]), .Ci(pp[06][10]), .S(fs[4]), .Co(fc[4]));
  fa fa5  (.A(pp[02][15]), .B(pp[03][14]), .Ci(pp[04][13]), .S(fs[5]), .Co(fc[5]));
  fa fa6  (.A(pp[05][12]), .B(pp[06][11]), .Ci(pp[07][10]), .S(fs[6]), .Co(fc[6]));
  fa fa7  (.A(pp[03][15]), .B(pp[04][14]), .Ci(pp[05][13]), .S(fs[7]), .Co(fc[7]));

  ha ha0  (.A(pp[00][13]), .B(pp[01][12]), .S(hs[0]), .C(hc[0]));
  ha ha1  (.A(pp[03][11]), .B(pp[04][10]), .S(hs[1]), .C(hc[1]));
  ha ha2  (.A(pp[06][09]), .B(pp[07][08]), .S(hs[2]), .C(hc[2]));
  ha ha3  (.A(pp[07][09]), .B(pp[08][08]), .S(hs[3]), .C(hc[3]));
  
  ////////////////////////////// RS2 16 -> 13 -> 9 /////////////////////////////
  // Adders : FA = 40; HA = 4;
  
  fa fa8  (.A(pp[00][10]), .B(pp[01][09]), .Ci(pp[02][08]), .S(fs[8]), .Co(fc[8]));
  fa fa9  (.A(pp[00][11]), .B(pp[01][10]), .Ci(pp[02][09]), .S(fs[9]), .Co(fc[9]));
  fa fa10 (.A(pp[03][08]), .B(pp[04][07]), .Ci(pp[05][06]), .S(fs[10]), .Co(fc[10]));
  fa fa11 (.A(pp[00][12]), .B(pp[01][11]), .Ci(pp[02][10]), .S(fs[11]), .Co(fc[11]));
  fa fa12 (.A(pp[03][09]), .B(pp[04][08]), .Ci(pp[05][07]), .S(fs[12]), .Co(fc[12]));
  fa fa13 (.A(pp[06][06]), .B(pp[07][05]), .Ci(pp[08][04]), .S(fs[13]), .Co(fc[13]));
  fa fa14 (.A(hs[0]), .B(pp[02][11]), .Ci(pp[03][10]), .S(fs[14]), .Co(fc[14]));
  fa fa15 (.A(pp[04][09]), .B(pp[05][08]), .Ci(pp[06][07]), .S(fs[15]), .Co(fc[15]));
  fa fa16 (.A(pp[07][06]), .B(pp[08][05]), .Ci(pp[09][04]), .S(fs[16]), .Co(fc[16]));
  fa fa17 (.A(pp[10][03]), .B(pp[11][02]), .Ci(pp[12][01]), .S(fs[17]), .Co(fc[17]));
  fa fa18 (.A(hc[0]), .B(fs[0]), .Ci(hs[1]), .S(fs[18]), .Co(fc[18]));
  fa fa19 (.A(pp[05][09]), .B(pp[06][08]), .Ci(pp[07][07]), .S(fs[19]), .Co(fc[19]));
  fa fa20 (.A(pp[08][06]), .B(pp[09][05]), .Ci(pp[10][04]), .S(fs[20]), .Co(fc[20]));
  fa fa21 (.A(pp[11][03]), .B(pp[12][02]), .Ci(pp[13][01]), .S(fs[21]), .Co(fc[21]));
  fa fa22 (.A(fc[0]), .B(hc[1]), .Ci(fs[1]), .S(fs[22]), .Co(fc[22]));
  fa fa23 (.A(fs[2]), .B(hs[2]), .Ci(pp[08][07]), .S(fs[23]), .Co(fc[23]));
  fa fa24 (.A(pp[09][06]), .B(pp[10][05]), .Ci(pp[11][04]), .S(fs[24]), .Co(fc[24]));
  fa fa25 (.A(pp[12][03]), .B(pp[13][02]), .Ci(pp[14][01]), .S(fs[25]), .Co(fc[25]));
  fa fa26 (.A(fc[1]), .B(fc[2]), .Ci(hc[2]), .S(fs[26]), .Co(fc[26]));
  fa fa27 (.A(fs[3]), .B(fs[4]), .Ci(hs[3]), .S(fs[27]), .Co(fc[27]));
  fa fa28 (.A(pp[09][07]), .B(pp[10][06]), .Ci(pp[11][05]), .S(fs[28]), .Co(fc[28]));
  fa fa29 (.A(pp[12][04]), .B(pp[13][03]), .Ci(pp[14][02]), .S(fs[29]), .Co(fc[29]));
  fa fa30 (.A(fc[3]), .B(fc[4]), .Ci(hc[3]), .S(fs[30]), .Co(fc[30]));
  fa fa31 (.A(fs[5]), .B(fs[6]), .Ci(pp[08][09]), .S(fs[31]), .Co(fc[31]));
  fa fa32 (.A(pp[09][08]), .B(pp[10][07]), .Ci(pp[11][06]), .S(fs[32]), .Co(fc[32]));
  fa fa33 (.A(pp[12][05]), .B(pp[13][04]), .Ci(pp[14][03]), .S(fs[33]), .Co(fc[33]));
  fa fa34 (.A(fc[5]), .B(fc[6]), .Ci(fs[7]), .S(fs[34]), .Co(fc[34]));
  fa fa35 (.A(pp[06][12]), .B(pp[07][11]), .Ci(pp[08][10]), .S(fs[35]), .Co(fc[35]));
  fa fa36 (.A(pp[09][09]), .B(pp[10][08]), .Ci(pp[11][07]), .S(fs[36]), .Co(fc[36]));
  fa fa37 (.A(pp[12][06]), .B(pp[13][05]), .Ci(pp[14][04]), .S(fs[37]), .Co(fc[37]));
  fa fa38 (.A(fc[7]), .B(pp[04][15]), .Ci(pp[05][14]), .S(fs[38]), .Co(fc[38]));
  fa fa39 (.A(pp[06][13]), .B(pp[07][12]), .Ci(pp[08][11]), .S(fs[39]), .Co(fc[39]));
  fa fa40 (.A(pp[09][10]), .B(pp[10][09]), .Ci(pp[11][08]), .S(fs[40]), .Co(fc[40]));
  fa fa41 (.A(pp[12][07]), .B(pp[13][06]), .Ci(pp[14][05]), .S(fs[41]), .Co(fc[41]));
  fa fa42 (.A(pp[05][15]), .B(pp[06][14]), .Ci(pp[07][13]), .S(fs[42]), .Co(fc[42]));
  fa fa43 (.A(pp[08][12]), .B(pp[09][11]), .Ci(pp[10][10]), .S(fs[43]), .Co(fc[43]));
  fa fa44 (.A(pp[11][09]), .B(pp[12][08]), .Ci(pp[13][07]), .S(fs[44]), .Co(fc[44]));
  fa fa45 (.A(pp[06][15]), .B(pp[07][14]), .Ci(pp[08][13]), .S(fs[45]), .Co(fc[45]));
  fa fa46 (.A(pp[09][12]), .B(pp[10][11]), .Ci(pp[11][10]), .S(fs[46]), .Co(fc[46]));
  fa fa47 (.A(pp[07][15]), .B(pp[08][14]), .Ci(pp[09][13]), .S(fs[47]), .Co(fc[47]));
  
  ha ha4  (.A(pp[00][09]), .B(pp[01][08]), .S(hs[4]), .C(hc[4]));
  ha ha5  (.A(pp[03][07]), .B(pp[04][06]), .S(hs[5]), .C(hc[5]));
  ha ha6  (.A(pp[06][05]), .B(pp[07][04]), .S(hs[6]), .C(hc[6]));
  ha ha7  (.A(pp[09][03]), .B(pp[10][02]), .S(hs[7]), .C(hc[7]));
  
  ////////////////////////////// RS3 16 -> 13 -> 9 -> 6/////////////////////////
  // Adders: FA = 51; HA = 3
  fa fa48 (.A(pp[00][07]), .B(pp[01][06]), .Ci(pp[02][05]), .S(fs[48]), .Co(fc[48]));
  fa fa49 (.A(pp[00][08]), .B(pp[01][07]), .Ci(pp[02][06]), .S(fs[49]), .Co(fc[49]));
  fa fa50 (.A(pp[03][05]), .B(pp[04][04]), .Ci(pp[05][03]), .S(fs[50]), .Co(fc[50]));
  fa fa51 (.A(hs[4]), .B(pp[02][07]), .Ci(pp[03][06]), .S(fs[51]), .Co(fc[51]));
  fa fa52 (.A(pp[04][05]), .B(pp[05][04]), .Ci(pp[06][03]), .S(fs[52]), .Co(fc[52]));
  fa fa53 (.A(pp[07][02]), .B(pp[08][01]), .Ci(pp[09][00]), .S(fs[53]), .Co(fc[53]));
  fa fa54 (.A(hc[4]), .B(fs[8]), .Ci(hs[5]), .S(fs[54]), .Co(fc[54]));
  fa fa55 (.A(pp[05][05]), .B(pp[06][04]), .Ci(pp[07][03]), .S(fs[55]), .Co(fc[55]));
  fa fa56 (.A(pp[08][02]), .B(pp[09][01]), .Ci(pp[10][00]), .S(fs[56]), .Co(fc[56]));
  fa fa57 (.A(fc[8]), .B(hc[5]), .Ci(fs[9]), .S(fs[57]), .Co(fc[57]));
  fa fa58 (.A(fs[10]), .B(hs[6]), .Ci(pp[08][03]), .S(fs[58]), .Co(fc[58]));
  fa fa59 (.A(pp[09][02]), .B(pp[10][01]), .Ci(pp[11][00]), .S(fs[59]), .Co(fc[59]));
  fa fa60 (.A(fc[9]), .B(fc[10]), .Ci(hc[6]), .S(fs[60]), .Co(fc[60]));
  fa fa61 (.A(fs[11]), .B(fs[12]), .Ci(fs[13]), .S(fs[61]), .Co(fc[61]));
  fa fa62 (.A(hs[7]), .B(pp[11][01]), .Ci(pp[12][00]), .S(fs[62]), .Co(fc[62]));
  fa fa63 (.A(fc[11]), .B(fc[12]), .Ci(fc[13]), .S(fs[63]), .Co(fc[63]));
  fa fa64 (.A(hc[7]), .B(fs[14]), .Ci(fs[15]), .S(fs[64]), .Co(fc[64]));
  fa fa65 (.A(fs[16]), .B(fs[17]), .Ci(pp[13][00]), .S(fs[65]), .Co(fc[65]));
  fa fa66 (.A(fc[14]), .B(fc[15]), .Ci(fc[16]), .S(fs[66]), .Co(fc[66]));
  fa fa67 (.A(fc[17]), .B(fs[18]), .Ci(fs[19]), .S(fs[67]), .Co(fc[67]));
  fa fa68 (.A(fs[20]), .B(fs[21]), .Ci(pp[14][00]), .S(fs[68]), .Co(fc[68]));
  fa fa69 (.A(fc[18]), .B(fc[19]), .Ci(fc[20]), .S(fs[69]), .Co(fc[69]));
  fa fa70 (.A(fc[21]), .B(fs[22]), .Ci(fs[23]), .S(fs[70]), .Co(fc[70]));
  fa fa71 (.A(fs[24]), .B(fs[25]), .Ci(pp[15][00]), .S(fs[71]), .Co(fc[71]));
  fa fa72 (.A(fc[22]), .B(fc[23]), .Ci(fc[24]), .S(fs[72]), .Co(fc[72]));
  fa fa73 (.A(fc[25]), .B(fs[26]), .Ci(fs[27]), .S(fs[73]), .Co(fc[73]));
  fa fa74 (.A(fs[28]), .B(fs[29]), .Ci(pp[15][01]), .S(fs[74]), .Co(fc[74]));
  fa fa75 (.A(fc[26]), .B(fc[27]), .Ci(fc[28]), .S(fs[75]), .Co(fc[75]));
  fa fa76 (.A(fc[29]), .B(fs[30]), .Ci(fs[31]), .S(fs[76]), .Co(fc[76]));
  fa fa77 (.A(fs[32]), .B(fs[33]), .Ci(pp[15][02]), .S(fs[77]), .Co(fc[77]));
  fa fa78 (.A(fc[30]), .B(fc[31]), .Ci(fc[32]), .S(fs[78]), .Co(fc[78]));
  fa fa79 (.A(fc[33]), .B(fs[34]), .Ci(fs[35]), .S(fs[79]), .Co(fc[79]));
  fa fa80 (.A(fs[36]), .B(fs[37]), .Ci(pp[15][03]), .S(fs[80]), .Co(fc[80]));
  fa fa81 (.A(fc[34]), .B(fc[35]), .Ci(fc[36]), .S(fs[81]), .Co(fc[81]));
  fa fa82 (.A(fc[37]), .B(fs[38]), .Ci(fs[39]), .S(fs[82]), .Co(fc[82]));
  fa fa83 (.A(fs[40]), .B(fs[41]), .Ci(pp[15][04]), .S(fs[83]), .Co(fc[83]));
  fa fa84 (.A(fc[38]), .B(fc[39]), .Ci(fc[40]), .S(fs[84]), .Co(fc[84]));
  fa fa85 (.A(fc[41]), .B(fs[42]), .Ci(fs[43]), .S(fs[85]), .Co(fc[85]));
  fa fa86 (.A(fs[44]), .B(pp[14][06]), .Ci(pp[15][05]), .S(fs[86]), .Co(fc[86]));
  fa fa87 (.A(fc[42]), .B(fc[43]), .Ci(fc[44]), .S(fs[87]), .Co(fc[87]));
  fa fa88 (.A(fs[45]), .B(fs[46]), .Ci(pp[12][09]), .S(fs[88]), .Co(fc[88]));
  fa fa89 (.A(pp[13][08]), .B(pp[14][07]), .Ci(pp[15][06]), .S(fs[89]), .Co(fc[89]));
  fa fa90 (.A(fc[45]), .B(fc[46]), .Ci(fs[47]), .S(fs[90]), .Co(fc[90]));
  fa fa91 (.A(pp[10][12]), .B(pp[11][11]), .Ci(pp[12][10]), .S(fs[91]), .Co(fc[91]));
  fa fa92 (.A(pp[13][09]), .B(pp[14][08]), .Ci(pp[15][07]), .S(fs[92]), .Co(fc[92]));
  fa fa93 (.A(fc[47]), .B(pp[08][15]), .Ci(pp[09][14]), .S(fs[93]), .Co(fc[93]));
  fa fa94 (.A(pp[10][13]), .B(pp[11][12]), .Ci(pp[12][11]), .S(fs[94]), .Co(fc[94]));
  fa fa95 (.A(pp[13][10]), .B(pp[14][09]), .Ci(pp[15][08]), .S(fs[95]), .Co(fc[95]));
  fa fa96 (.A(pp[09][15]), .B(pp[10][14]), .Ci(pp[11][13]), .S(fs[96]), .Co(fc[96]));
  fa fa97 (.A(pp[12][12]), .B(pp[13][11]), .Ci(pp[14][10]), .S(fs[97]), .Co(fc[97]));
  fa fa98 (.A(pp[10][15]), .B(pp[11][14]), .Ci(pp[12][13]), .S(fs[98]), .Co(fc[98]));
  
  ha ha8  (.A(pp[00][06]), .B(pp[01][05]), .S(hs[ 8]), .C(hc[8]));
  ha ha9  (.A(pp[03][04]), .B(pp[04][03]), .S(hs[ 9]), .C(hc[9]));
  ha ha10 (.A(pp[06][02]), .B(pp[07][01]), .S(hs[10]), .C(hc[10]));
  
  ////////////////////////////// RS4 16 -> 13 -> 9 -> 6 -> 4////////////////////
  //Adders: FA = 44; HA = 2
  
  fa fa99  (.A(pp[00][05]), .B(pp[01][04]), .Ci(pp[02][03]), .S(fs[99]), .Co(fc[99]));
  fa fa100 (.A(hs[8]), .B(pp[02][04]), .Ci(pp[03][03]), .S(fs[100]), .Co(fc[100]));
  fa fa101 (.A(pp[04][02]), .B(pp[05][01]), .Ci(pp[06][00]), .S(fs[101]), .Co(fc[101]));
  fa fa102 (.A(hc[8]), .B(fs[48]), .Ci(hs[9]), .S(fs[102]), .Co(fc[102]));
  fa fa103 (.A(pp[05][02]), .B(pp[06][01]), .Ci(pp[07][00]), .S(fs[103]), .Co(fc[103]));
  fa fa104 (.A(fc[48]), .B(hc[9]), .Ci(fs[49]), .S(fs[104]), .Co(fc[104]));
  fa fa105 (.A(fs[50]), .B(hs[10]), .Ci(pp[08][00]), .S(fs[105]), .Co(fc[105]));
  fa fa106 (.A(fc[49]), .B(fc[50]), .Ci(hc[10]), .S(fs[106]), .Co(fc[106]));
  fa fa107 (.A(fs[51]), .B(fs[52]), .Ci(fs[53]), .S(fs[107]), .Co(fc[107]));
  fa fa108 (.A(fc[51]), .B(fc[52]), .Ci(fc[53]), .S(fs[108]), .Co(fc[108]));
  fa fa109 (.A(fs[54]), .B(fs[55]), .Ci(fs[56]), .S(fs[109]), .Co(fc[109]));
  fa fa110 (.A(fc[54]), .B(fc[55]), .Ci(fc[56]), .S(fs[110]), .Co(fc[110]));
  fa fa111 (.A(fs[57]), .B(fs[58]), .Ci(fs[59]), .S(fs[111]), .Co(fc[111]));
  fa fa112 (.A(fc[57]), .B(fc[58]), .Ci(fc[59]), .S(fs[112]), .Co(fc[112]));
  fa fa113 (.A(fs[60]), .B(fs[61]), .Ci(fs[62]), .S(fs[113]), .Co(fc[113]));
  fa fa114 (.A(fc[60]), .B(fc[61]), .Ci(fc[62]), .S(fs[114]), .Co(fc[114]));
  fa fa115 (.A(fs[63]), .B(fs[64]), .Ci(fs[65]), .S(fs[115]), .Co(fc[115]));
  fa fa116 (.A(fc[63]), .B(fc[64]), .Ci(fc[65]), .S(fs[116]), .Co(fc[116]));
  fa fa117 (.A(fs[66]), .B(fs[67]), .Ci(fs[68]), .S(fs[117]), .Co(fc[117]));
  fa fa118 (.A(fc[66]), .B(fc[67]), .Ci(fc[68]), .S(fs[118]), .Co(fc[118]));
  fa fa119 (.A(fs[69]), .B(fs[70]), .Ci(fs[71]), .S(fs[119]), .Co(fc[119]));
  fa fa120 (.A(fc[69]), .B(fc[70]), .Ci(fc[71]), .S(fs[120]), .Co(fc[120]));
  fa fa121 (.A(fs[72]), .B(fs[73]), .Ci(fs[74]), .S(fs[121]), .Co(fc[121]));
  fa fa122 (.A(fc[72]), .B(fc[73]), .Ci(fc[74]), .S(fs[122]), .Co(fc[122]));
  fa fa123 (.A(fs[75]), .B(fs[76]), .Ci(fs[77]), .S(fs[123]), .Co(fc[123]));
  fa fa124 (.A(fc[75]), .B(fc[76]), .Ci(fc[77]), .S(fs[124]), .Co(fc[124]));
  fa fa125 (.A(fs[78]), .B(fs[79]), .Ci(fs[80]), .S(fs[125]), .Co(fc[125]));
  fa fa126 (.A(fc[78]), .B(fc[79]), .Ci(fc[80]), .S(fs[126]), .Co(fc[126]));
  fa fa127 (.A(fs[81]), .B(fs[82]), .Ci(fs[83]), .S(fs[127]), .Co(fc[127]));
  fa fa128 (.A(fc[81]), .B(fc[82]), .Ci(fc[83]), .S(fs[128]), .Co(fc[128]));
  fa fa129 (.A(fs[84]), .B(fs[85]), .Ci(fs[86]), .S(fs[129]), .Co(fc[129]));
  fa fa130 (.A(fc[84]), .B(fc[85]), .Ci(fc[86]), .S(fs[130]), .Co(fc[130]));
  fa fa131 (.A(fs[87]), .B(fs[88]), .Ci(fs[89]), .S(fs[131]), .Co(fc[131]));
  fa fa132 (.A(fc[87]), .B(fc[88]), .Ci(fc[89]), .S(fs[132]), .Co(fc[132]));
  fa fa133 (.A(fs[90]), .B(fs[91]), .Ci(fs[92]), .S(fs[133]), .Co(fc[133]));
  fa fa134 (.A(fc[90]), .B(fc[91]), .Ci(fc[92]), .S(fs[134]), .Co(fc[134]));
  fa fa135 (.A(fs[93]), .B(fs[94]), .Ci(fs[95]), .S(fs[135]), .Co(fc[135]));
  fa fa136 (.A(fc[93]), .B(fc[94]), .Ci(fc[95]), .S(fs[136]), .Co(fc[136]));
  fa fa137 (.A(fs[96]), .B(fs[97]), .Ci(pp[15][09]), .S(fs[137]), .Co(fc[137]));
  fa fa138 (.A(fc[96]), .B(fc[97]), .Ci(fs[98]), .S(fs[138]), .Co(fc[138]));
  fa fa139 (.A(pp[13][12]), .B(pp[14][11]), .Ci(pp[15][10]), .S(fs[139]), .Co(fc[139]));
  fa fa140 (.A(fc[98]), .B(pp[11][15]), .Ci(pp[12][14]), .S(fs[140]), .Co(fc[140]));
  fa fa141 (.A(pp[13][13]), .B(pp[14][12]), .Ci(pp[15][11]), .S(fs[141]), .Co(fc[141]));
  fa fa142 (.A(pp[12][15]), .B(pp[13][14]), .Ci(pp[14][13]), .S(fs[142]), .Co(fc[142]));
  
   ha ha11   (.A(pp[00][04]), .B(pp[01][03]), .S(hs[11]), .C(hc[11]));
   ha ha12   (.A(pp[03][02]), .B(pp[04][01]), .S(hs[12]), .C(hc[12]));
    
  ///////////////////////////// RS5 16 -> 13 -> 9 -> 6 -> 4 -> 3////////////////
 
 // Adders: FA = 25; HA = 1
 
 fa fa143 (.A(hs[11]), .B(pp[02][02]), .Ci(pp[03][01]), .S(fs[143]), .Co(fc[143]));
 fa fa144 (.A(hc[11]), .B(fs[99]), .Ci(hs[12]), .S(fs[144]), .Co(fc[144]));
 fa fa145 (.A(fc[99]), .B(hc[12]), .Ci(fs[100]), .S(fs[145]), .Co(fc[145]));
 fa fa146 (.A(fc[100]), .B(fc[101]), .Ci(fs[102]), .S(fs[146]), .Co(fc[146]));
 fa fa147 (.A(fc[102]), .B(fc[103]), .Ci(fs[104]), .S(fs[147]), .Co(fc[147]));
 fa fa148 (.A(fc[104]), .B(fc[105]), .Ci(fs[106]), .S(fs[148]), .Co(fc[148]));
 fa fa149 (.A(fc[106]), .B(fc[107]), .Ci(fs[108]), .S(fs[149]), .Co(fc[149]));
 fa fa150 (.A(fc[108]), .B(fc[109]), .Ci(fs[110]), .S(fs[150]), .Co(fc[150]));
 fa fa151 (.A(fc[110]), .B(fc[111]), .Ci(fs[112]), .S(fs[151]), .Co(fc[151]));
 fa fa152 (.A(fc[112]), .B(fc[113]), .Ci(fs[114]), .S(fs[152]), .Co(fc[152]));
 fa fa153 (.A(fc[114]), .B(fc[115]), .Ci(fs[116]), .S(fs[153]), .Co(fc[153]));
 fa fa154 (.A(fc[116]), .B(fc[117]), .Ci(fs[118]), .S(fs[154]), .Co(fc[154]));
 fa fa155 (.A(fc[118]), .B(fc[119]), .Ci(fs[120]), .S(fs[155]), .Co(fc[155]));
 fa fa156 (.A(fc[120]), .B(fc[121]), .Ci(fs[122]), .S(fs[156]), .Co(fc[156]));
 fa fa157 (.A(fc[122]), .B(fc[123]), .Ci(fs[124]), .S(fs[157]), .Co(fc[157]));
 fa fa158 (.A(fc[124]), .B(fc[125]), .Ci(fs[126]), .S(fs[158]), .Co(fc[158]));
 fa fa159 (.A(fc[126]), .B(fc[127]), .Ci(fs[128]), .S(fs[159]), .Co(fc[159]));
 fa fa160 (.A(fc[128]), .B(fc[129]), .Ci(fs[130]), .S(fs[160]), .Co(fc[160]));
 fa fa161 (.A(fc[130]), .B(fc[131]), .Ci(fs[132]), .S(fs[161]), .Co(fc[161]));
 fa fa162 (.A(fc[132]), .B(fc[133]), .Ci(fs[134]), .S(fs[162]), .Co(fc[162]));
 fa fa163 (.A(fc[134]), .B(fc[135]), .Ci(fs[136]), .S(fs[163]), .Co(fc[163]));
 fa fa164 (.A(fc[136]), .B(fc[137]), .Ci(fs[138]), .S(fs[164]), .Co(fc[164]));
 fa fa165 (.A(fc[138]), .B(fc[139]), .Ci(fs[140]), .S(fs[165]), .Co(fc[165]));
 fa fa166 (.A(fc[140]), .B(fc[141]), .Ci(fs[142]), .S(fs[166]), .Co(fc[166]));
 fa fa167 (.A(fc[142]), .B(pp[13][15]), .Ci(pp[14][14]), .S(fs[167]), .Co(fc[167]));
 
 ha ha13  (.A(pp[00][03]), .B(pp[01][02]), .S(hs[13]), .C(hc[13]));
 
  ///////////////////////////// RS6 16 -> 13 -> 9 -> 6 -> 4 -> 3 -> 2///////////
  // Adders: FA = 27; HA = 1
  
   fa fa168 (.A(hs[13]), .B(pp[02][01]), .Ci(pp[03][00]), .S(to_FA[1][3]), .Co(to_FA[0][4]));
   fa fa169 (.A(hc[13]), .B(fs[143]), .Ci(pp[04][00]), .S(to_FA[1][4]), .Co(to_FA[0][5]));
   fa fa170 (.A(fc[143]), .B(fs[144]), .Ci(pp[05][00]), .S(to_FA[1][5]), .Co(to_FA[0][6]));
   fa fa171 (.A(fc[144]), .B(fs[145]), .Ci(fs[101]), .S(to_FA[1][6]),  .Co(to_FA[0][7]));
   fa fa172 (.A(fc[145]), .B(fs[146]), .Ci(fs[103]), .S(to_FA[1][7]),  .Co(to_FA[0][8]));
   fa fa173 (.A(fc[146]), .B(fs[147]), .Ci(fs[105]), .S(to_FA[1][8]),  .Co(to_FA[0][9]));
   fa fa174 (.A(fc[147]), .B(fs[148]), .Ci(fs[107]), .S(to_FA[1][9]),  .Co(to_FA[0][10]));
   fa fa175 (.A(fc[148]), .B(fs[149]), .Ci(fs[109]), .S(to_FA[1][10]), .Co(to_FA[0][11]));
   fa fa176 (.A(fc[149]), .B(fs[150]), .Ci(fs[111]), .S(to_FA[1][11]), .Co(to_FA[0][12]));
   fa fa177 (.A(fc[150]), .B(fs[151]), .Ci(fs[113]), .S(to_FA[1][12]), .Co(to_FA[0][13]));
   fa fa178 (.A(fc[151]), .B(fs[152]), .Ci(fs[115]), .S(to_FA[1][13]), .Co(to_FA[0][14]));
   fa fa179 (.A(fc[152]), .B(fs[153]), .Ci(fs[117]), .S(to_FA[1][14]), .Co(to_FA[0][15]));
   fa fa180 (.A(fc[153]), .B(fs[154]), .Ci(fs[119]), .S(to_FA[1][15]), .Co(to_FA[0][16]));
   fa fa181 (.A(fc[154]), .B(fs[155]), .Ci(fs[121]), .S(to_FA[1][16]), .Co(to_FA[0][17]));
   fa fa182 (.A(fc[155]), .B(fs[156]), .Ci(fs[123]), .S(to_FA[1][17]), .Co(to_FA[0][18]));
   fa fa183 (.A(fc[156]), .B(fs[157]), .Ci(fs[125]), .S(to_FA[1][18]), .Co(to_FA[0][19]));
   fa fa184 (.A(fc[157]), .B(fs[158]), .Ci(fs[127]), .S(to_FA[1][19]), .Co(to_FA[0][20]));
   fa fa185 (.A(fc[158]), .B(fs[159]), .Ci(fs[129]), .S(to_FA[1][20]), .Co(to_FA[0][21]));
   fa fa186 (.A(fc[159]), .B(fs[160]), .Ci(fs[131]), .S(to_FA[1][21]), .Co(to_FA[0][22]));
   fa fa187 (.A(fc[160]), .B(fs[161]), .Ci(fs[133]), .S(to_FA[1][22]), .Co(to_FA[0][23]));
   fa fa188 (.A(fc[161]), .B(fs[162]), .Ci(fs[135]), .S(to_FA[1][23]), .Co(to_FA[0][24]));
   fa fa189 (.A(fc[162]), .B(fs[163]), .Ci(fs[137]), .S(to_FA[1][24]), .Co(to_FA[0][25]));
   fa fa190 (.A(fc[163]), .B(fs[164]), .Ci(fs[139]), .S(to_FA[1][25]), .Co(to_FA[0][26]));
   fa fa191 (.A(fc[164]), .B(fs[165]), .Ci(fs[141]), .S(to_FA[1][26]), .Co(to_FA[0][27]));
   fa fa192 (.A(fc[165]), .B(fs[166]), .Ci(pp[15][12]), .S(to_FA[1][27]), .Co(to_FA[0][28]));
   fa fa193 (.A(fc[166]), .B(fs[167]), .Ci(pp[15][13]), .S(to_FA[1][28]), .Co(to_FA[0][29]));
   fa fa194 (.A(fc[167]), .B(pp[14][15]), .Ci(pp[15][14]), .S(to_FA[1][29]), .Co(to_FA[0][30]));
   
   ha ha14  (.A(pp[00][02]), .B(pp[01][01]), .S(to_FA[0][2]), .C(to_FA[0][3]));
  
  //mapping outputs
  assign to_FA[0][0] = pp[00][00];
  assign to_FA[1][0] = 1'b0;
  
  assign to_FA[0][1] = pp[00][01];
  assign to_FA[1][1] = pp[01][00];
  
  assign to_FA[1][2] = pp[02][00];
  
  assign to_FA[1][30] = pp[15][15]; 
  
  assign to_FA[0][31] = 1'b0;
  assign to_FA[1][31] = 1'b0; 
  
endmodule


////////////////////////////////////// 16 bit approximate multipliers processing blocks //////

module processing_block_16_1step(
input p[15:0][15:0],
output [30:0]out1,
output [30:0]out2);
      
    ////////////////////////////////////////// PP REDUCTION STEP ONE   ////////////////////////  
    wire r1[30:0][11:0] ; // outputs of first reduction
    
    assign r1[0][0] = p[0][0];                                                 // column 0
    assign r1[1][0] = p[1][0]; assign r1[1][1] = p[0][1];                       // column 1
    compressor3_2 c1   (.p({p[2][0]  ,p[1][1]  ,p[0][2]}),                                                                                                                    .w({r1[2][0] ,r1[2][1]}));                                                // column 2
    compressor4_2 c2   (.p({p[3][0]  ,p[2][1]  ,p[1][2] ,p[0][3]}),                                                                                                           .w({r1[3][0] ,r1[3][1]}));                                              // column 3
    compressor5_3 c3   (.p({p[4][0]  ,p[3][1]  ,p[2][2] ,p[1][3] ,p[0][4]}),                                                                                                  .w({r1[4][0] ,r1[4][1] ,r1[4][2]}));                                      // column 4
    compressor6_3 c4   (.p({p[5][0]  ,p[4][1]  ,p[3][2] ,p[2][3] ,p[1][4]  ,p[0][5]}),                                                                                        .w({r1[5][0] ,r1[5][1] ,r1[5][2]}));                                    // column 5
    compressor7_4 c5   (.p({p[6][0]  ,p[5][1]  ,p[4][2] ,p[3][3] ,p[2][4]  ,p[1][5] ,p[0][6]}),                                                                               .w({r1[6][0] ,r1[6][1] ,r1[6][2] ,r1[6][3]}));                               // column 6
    compressor8_4 c6   (.p({p[7][0]  ,p[6][1]  ,p[5][2] ,p[4][3] ,p[3][4]  ,p[2][5] ,p[1][6],p[0][7]}),                                                                       .w({r1[7][0] ,r1[7][1] ,r1[7][2] ,r1[7][3]}));                                // column 7
    compressor9_5 c7   (.p({p[8][0]  ,p[7][1]  ,p[6][2] ,p[5][3] ,p[4][4]  ,p[3][5] ,p[2][6],p[1][7],p[0][8]}),                                                               .w({r1[8][0] ,r1[8][1] ,r1[8][2] ,r1[8][3] ,r1[8][4]}));                       // column 8
    compressor10_5 c8  (.p({p[9][0]  ,p[8][1]  ,p[7][2] ,p[6][3] ,p[5][4]  ,p[4][5] ,p[3][6],p[2][7],p[1][8],p[0][9]}),                                                       .w({r1[9][0] ,r1[9][1] ,r1[9][2] ,r1[9][3] ,r1[9][4]}));                         // column 9
    compressor11_6 c9  (.p({p[10][0] ,p[9][1]  ,p[8][2] ,p[7][3] ,p[6][4]  ,p[5][5] ,p[4][6],p[3][7],p[2][8],p[1][9],p[0][10]}),                                              .w({r1[10][0],r1[10][1],r1[10][2],r1[10][3],r1[10][4],r1[10][5]}));              // column 10
    compressor12_6 c10 (.p({p[11][0] ,p[10][1] ,p[9][2] ,p[8][3] ,p[7][4]  ,p[6][5] ,p[5][6],p[4][7],p[3][8],p[2][9],p[1][10],p[0][11]}),                                     .w({r1[11][0],r1[11][1],r1[11][2],r1[11][3],r1[11][4],r1[11][5]}));              // column 11
    compressor13_7 c11 (.p({p[12][0] ,p[11][1] ,p[10][2],p[9][3] ,p[8][4]  ,p[7][5] ,p[6][6],p[5][7],p[4][8],p[3][9],p[2][10],p[1][11],p[0][12]}),                            .w({r1[12][0],r1[12][1],r1[12][2],r1[12][3],r1[12][4],r1[12][5],r1[12][6]}));     // column 12
    compressor14_7 c12 (.p({p[13][0] ,p[12][1] ,p[11][2],p[10][3],p[9][4]  ,p[8][5] ,p[7][6],p[6][7],p[5][8],p[4][9],p[3][10],p[2][11],p[1][12],p[0][13]}),                   .w({r1[13][0],r1[13][1],r1[13][2],r1[13][3],r1[13][4],r1[13][5],r1[13][6]}));      // column 13
    compressor15_8 c13 (.p({p[14][0] ,p[13][1] ,p[12][2],p[11][3],p[10][4] ,p[9][5] ,p[8][6],p[7][7],p[6][8],p[5][9],p[4][10],p[3][11],p[2][12],p[1][13],p[0][14]}),          .w({r1[14][0],r1[14][1],r1[14][2],r1[14][3],r1[14][4],r1[14][5],r1[14][6],r1[14][7]})); // column 14
    compressor16_8 c14 (.p({p[15][0] ,p[14][1] ,p[13][2],p[12][3],p[11][4] ,p[10][5],p[9][6],p[8][7],p[7][8],p[6][9],p[5][10],p[4][11],p[3][12],p[2][13],p[1][14],p[0][15]}), .w({r1[15][0],r1[15][1],r1[15][2],r1[15][3],r1[15][4],r1[15][5],r1[15][6],r1[15][7]})); // column 15
    
    compressor14_7 c15 (.p({p[15][1] ,p[14][2] ,p[13][3],p[12][4],p[11][5]  ,p[10][6] ,p[9][7],p[8][8],p[7][9],p[6][10],p[5][11],p[4][12],p[3][13],p[2][14]}),                .w({r1[16][0],r1[16][1],r1[16][2],r1[16][3],r1[16][4],r1[16][5],r1[16][6]}));
    assign r1[16][7] = p[1][15];// column 16
    
    FA e1(.p({p[15][2],p[14][3],p[13][4]}), .w({r1[18][0],r1[17][0]})   );
    FA e2(.p({p[12][5],p[11][6],p[10][7]}), .w({r1[18][1],r1[17][1]})   );
    FA e3(.p({p[9][8],p[8][9],p[7][10]}), .w({r1[18][2],r1[17][2]})   ); 
    assign r1[17][3] = p[6][11];
    assign r1[17][4] = p[5][12];
    assign r1[17][5] = p[4][13];
    assign r1[17][6] = p[3][14];
    assign r1[17][7] = p[2][15];//column 17
    
    FA e4(.p({p[15][3],p[14][4],p[13][5]}), .w({r1[19][0],r1[18][3]})   );
    FA e5(.p({p[12][6],p[11][7],p[10][8]}), .w({r1[19][1],r1[18][4]})   );
    FA e6(.p({p[9][9],p[8][10],p[7][11]}), .w({r1[19][2],r1[18][5]})   ); 
    FA e7(.p({p[6][12],p[5][13],p[4][14]}), .w({r1[19][3],r1[18][6]})   );
    assign r1[18][7] = p[3][15]; //column 18
    
    FA e8(.p({p[15][4],p[14][5],p[13][6]}),  .w({r1[20][0],r1[19][4]})   );
    FA e9(.p({p[12][7],p[11][8],p[10][9]}),  .w({r1[20][1],r1[19][5]})   );
    FA e10(.p({p[9][10],p[8][11],p[7][12]}), .w({r1[20][2],r1[19][6]})   ); 
    FA e11(.p({p[6][13],p[5][14],p[4][15]}), .w({r1[20][3],r1[19][7]})   ); //column 19
    
    FA e12(.p({p[15][5],p[14][6],p[13][7]}),  .w({r1[21][0],r1[20][4]})   );
    FA e13(.p({p[12][8],p[11][9],p[10][10]}), .w({r1[21][1],r1[20][5]})   );
    FA e14(.p({p[9][11],p[8][12],p[7][13]}),  .w({r1[21][2],r1[20][6]})   );
    HA e15(.p({p[6][14],p[5][15]}),           .w({r1[21][3],r1[20][7]})   ); //column 20
    
    FA e16(.p({p[15][6],p[14][7],p[13][8]}),   .w({r1[22][0],r1[21][4]})   );
    FA e17(.p({p[12][9],p[11][10],p[10][11]}), .w({r1[22][1],r1[21][5]})   );
    FA e18(.p({p[9][12],p[8][13],p[7][14]}),   .w({r1[22][2],r1[21][6]})   );
    assign r1[21][7] = p[6][15]; //column 21
    
    FA e19(.p({p[15][7],p[14][8],p[13][9]}),    .w({r1[23][0],r1[22][3]})   );
    FA e20(.p({p[12][10],p[11][11],p[10][12]}), .w({r1[23][1],r1[22][4]})   ); 
    assign r1[22][5] = p[9][13];
    assign r1[22][6] = p[8][14];
    assign r1[22][7] = p[7][15]; //column 22
    
    FA e21(.p({p[15][8],p[14][9],p[13][10]}), .w({r1[24][0],r1[23][2]})   );
    assign r1[23][3] = p[12][11];
    assign r1[23][4] = p[11][12];
    assign r1[23][5] = p[10][13];
    assign r1[23][6] = p[9][14];
    assign r1[23][7] = p[8][15]; //column 23
    
    assign r1[24][1] = p[15][9];
    assign r1[24][2] = p[14][10];
    assign r1[24][3] = p[13][11];
    assign r1[24][4] = p[12][12];
    assign r1[24][5] = p[11][13];
    assign r1[24][6] = p[10][14];
    assign r1[24][7] = p[9][15]; //column 24
    
    assign r1[25][0] = p[15][10];
    assign r1[25][1] = p[14][11];
    assign r1[25][2] = p[13][12];
    assign r1[25][3] = p[12][13];
    assign r1[25][4] = p[11][14];
    assign r1[25][5] = p[10][15]; //column 25
    
    assign r1[26][0] = p[15][11];
    assign r1[26][1] = p[14][12];
    assign r1[26][2] = p[13][13];
    assign r1[26][3] = p[12][14];
    assign r1[26][4] = p[11][15]; //column 26
    
    assign r1[27][0] = p[15][12];
    assign r1[27][1] = p[14][13];
    assign r1[27][2] = p[13][14];
    assign r1[27][3] = p[12][15]; //column 27
    
    assign r1[28][0] = p[15][13];
    assign r1[28][1] = p[14][14];
    assign r1[28][2] = p[13][15]; //column 28
    
    assign r1[29][0] = p[15][14];
    assign r1[29][1] = p[14][15]; //column 29
   
    assign r1[30][0] = p[15][15]; //column 30
    
    
    ////////////////////////////////////////// exact adders one   ////////////////////////  
    wire r2[30:0][5:0] ; // outputs of first reduction
	
	assign r2[0][0] = r1[0][0]; // column 0
	
	assign r2[1][0] = r1[1][0];
	assign r2[1][1] = r1[1][1]; // column 1
	
	assign r2[2][0] = r1[2][0];
	assign r2[2][1] = r1[2][1]; // column 2
	
	assign r2[3][0] = r1[3][0];
	assign r2[3][1] = r1[3][1]; // column 3
	
	assign r2[4][1] = 1'b0;
	FA e22(.p({r1[4][0],r1[4][1],r1[4][2]}),    .w({r1[5][3],r2[4][0]})   ); // column 4
	
	assign r2[5][1] = r1[5][3];
	FA e23(.p({r1[5][0],r1[5][1],r1[5][2]}),    .w({r1[6][4],r2[5][0]})   ); // column 5
	
	FA e24(.p({r1[6][0],r1[6][1],r1[6][2]}),    .w({r1[7][4],r2[6][0]})   );
	HA e25(.p({r1[6][3],r1[6][4]}),             .w({r1[7][5],r2[6][1]})   ); // column 6
	
	FA e26(.p({r1[7][0],r1[7][1],r1[7][2]}),    .w({r1[8][5],r2[7][0]})   );
	FA e27(.p({r1[7][3],r1[7][4],r1[7][5]}),    .w({r1[8][6],r2[7][1]})   ); // column 7
	
	assign r2[8][2] = r1[8][6];
	FA e28(.p({r1[8][0],r1[8][1],r1[8][2]}),    .w({r1[9][5],r2[8][0]})   );
	FA e29(.p({r1[8][3],r1[8][4],r1[8][5]}),    .w({r1[9][6],r2[8][1]})   ); // column 8
	
	assign r2[9][2] = r1[9][6];
	FA e30(.p({r1[9][0],r1[9][1],r1[9][2]}),    .w({r1[10][6],r2[9][0]})   );
	FA e31(.p({r1[9][3],r1[9][4],r1[9][5]}),    .w({r1[10][7],r2[9][1]})   ); // column 9
	
	FA e32(.p({r1[10][0],r1[10][1],r1[10][2]}),    .w({r1[11][6],r2[10][0]})   );
	FA e33(.p({r1[10][3],r1[10][4],r1[10][5]}),    .w({r1[11][7],r2[10][1]})   );
	HA e34(.p({r1[10][6],r1[10][7]}),              .w({r1[11][8],r2[10][2]})   ); // column 10
	
	FA e35(.p({r1[11][0],r1[11][1],r1[11][2]}),    .w({r1[12][7],r2[11][0]})   );
	FA e36(.p({r1[11][3],r1[11][4],r1[11][5]}),    .w({r1[12][8],r2[11][1]})   );
	FA e37(.p({r1[11][6],r1[11][7],r1[11][8]}),    .w({r1[12][9],r2[11][2]})   ); // column 11
	
	assign r2[12][3] = r1[12][9];
	FA e38(.p({r1[12][0],r1[12][1],r1[12][2]}),    .w({r1[13][7],r2[12][0]})   );
	FA e39(.p({r1[12][3],r1[12][4],r1[12][5]}),    .w({r1[13][8],r2[12][1]})   );
	FA e40(.p({r1[12][6],r1[12][7],r1[12][8]}),    .w({r1[13][9],r2[12][2]})   ); // column 12
	
	assign r2[13][3] = r1[13][9];
	FA e41(.p({r1[13][0],r1[13][1],r1[13][2]}),    .w({r1[14][8 ],r2[13][0]})   );
	FA e42(.p({r1[13][3],r1[13][4],r1[13][5]}),    .w({r1[14][9 ],r2[13][1]})   );
	FA e43(.p({r1[13][6],r1[13][7],r1[13][8]}),    .w({r1[14][10],r2[13][2]})   ); // column 13
	
	FA e44(.p({r1[14][0],r1[14][1],r1[14][2]}),    .w({r1[15][8 ],r2[14][0]})   );
	FA e45(.p({r1[14][3],r1[14][4],r1[14][5]}),    .w({r1[15][9 ],r2[14][1]})   );
	FA e46(.p({r1[14][6],r1[14][7],r1[14][8]}),    .w({r1[15][10],r2[14][2]})   );
	HA e47(.p({r1[14][9],r1[14][10]}),             .w({r1[15][11],r2[14][3]})   ); // column 14
	
	FA e48(.p({r1[15][0],r1[15][1 ],r1[15][2 ]}),    .w({r1[16][8 ],r2[15][0]})   );
	FA e49(.p({r1[15][3],r1[15][4 ],r1[15][5 ]}),    .w({r1[16][9 ],r2[15][1]})   );
	FA e50(.p({r1[15][6],r1[15][7 ],r1[15][8 ]}),    .w({r1[16][10],r2[15][2]})   );
	FA e51(.p({r1[15][9],r1[15][10],r1[15][11]}),    .w({r1[16][11],r2[15][3]})   ); // column 15
	
	FA e52(.p({r1[16][0],r1[16][1 ],r1[16][2 ]}),    .w({r1[17][8 ],r2[16][0]})   );
	FA e53(.p({r1[16][3],r1[16][4 ],r1[16][5 ]}),    .w({r1[17][9 ],r2[16][1]})   );
	FA e54(.p({r1[16][6],r1[16][7 ],r1[16][8 ]}),    .w({r1[17][10],r2[16][2]})   );
	FA e55(.p({r1[16][9],r1[16][10],r1[16][11]}),    .w({r1[17][11],r2[16][3]})   ); // column 16
	
	FA e56(.p({r1[17][0],r1[17][1 ],r1[17][2 ]}),    .w({r1[18][8 ],r2[17][0]})   );
	FA e57(.p({r1[17][3],r1[17][4 ],r1[17][5 ]}),    .w({r1[18][9 ],r2[17][1]})   );
	FA e58(.p({r1[17][6],r1[17][7 ],r1[17][8 ]}),    .w({r1[18][10],r2[17][2]})   );
	FA e59(.p({r1[17][9],r1[17][10],r1[17][11]}),    .w({r1[18][11],r2[17][3]})   ); // column 17
	
	FA e60(.p({r1[18][0],r1[18][1 ],r1[18][2 ]}),    .w({r1[19][8 ],r2[18][0]})   );
	FA e61(.p({r1[18][3],r1[18][4 ],r1[18][5 ]}),    .w({r1[19][9 ],r2[18][1]})   );
	FA e62(.p({r1[18][6],r1[18][7 ],r1[18][8 ]}),    .w({r1[19][10],r2[18][2]})   );
	FA e63(.p({r1[18][9],r1[18][10],r1[18][11]}),    .w({r1[19][11],r2[18][3]})   ); // column 18
	
	FA e64(.p({r1[19][0],r1[19][1 ],r1[19][2 ]}),    .w({r1[20][8 ],r2[19][0]})   );
	FA e65(.p({r1[19][3],r1[19][4 ],r1[19][5 ]}),    .w({r1[20][9 ],r2[19][1]})   );
	FA e66(.p({r1[19][6],r1[19][7 ],r1[19][8 ]}),    .w({r1[20][10],r2[19][2]})   );
	FA e67(.p({r1[19][9],r1[19][10],r1[19][11]}),    .w({r1[20][11],r2[19][3]})   ); // column 19
	
	FA e68(.p({r1[20][0],r1[20][1 ],r1[20][2 ]}),    .w({r1[21][8 ],r2[20][0]})   );
	FA e69(.p({r1[20][3],r1[20][4 ],r1[20][5 ]}),    .w({r1[21][9 ],r2[20][1]})   );
	FA e70(.p({r1[20][6],r1[20][7 ],r1[20][8 ]}),    .w({r1[21][10],r2[20][2]})   );
	FA e71(.p({r1[20][9],r1[20][10],r1[20][11]}),    .w({r1[21][11],r2[20][3]})   ); // column 20
	
	FA e72(.p({r1[21][0],r1[21][1 ],r1[21][2 ]}),    .w({r1[22][8 ],r2[21][0]})   );
	FA e73(.p({r1[21][3],r1[21][4 ],r1[21][5 ]}),    .w({r1[22][9 ],r2[21][1]})   );
	FA e74(.p({r1[21][6],r1[21][7 ],r1[21][8 ]}),    .w({r1[22][10],r2[21][2]})   );
	FA e75(.p({r1[21][9],r1[21][10],r1[21][11]}),    .w({r1[22][11],r2[21][3]})   ); // column 21
	
	FA e76(.p({r1[22][0],r1[22][1 ],r1[22][2 ]}),    .w({r1[23][8 ],r2[22][0]})   );
	FA e77(.p({r1[22][3],r1[22][4 ],r1[22][5 ]}),    .w({r1[23][9 ],r2[22][1]})   );
	FA e78(.p({r1[22][6],r1[22][7 ],r1[22][8 ]}),    .w({r1[23][10],r2[22][2]})   );
	FA e79(.p({r1[22][9],r1[22][10],r1[22][11]}),    .w({r1[23][11],r2[22][3]})   ); // column 22
	
	FA e80(.p({r1[23][0],r1[23][1 ],r1[23][2 ]}),    .w({r1[24][8 ],r2[23][0]})   );
	FA e81(.p({r1[23][3],r1[23][4 ],r1[23][5 ]}),    .w({r1[24][9 ],r2[23][1]})   );
	FA e82(.p({r1[23][6],r1[23][7 ],r1[23][8 ]}),    .w({r1[24][10],r2[23][2]})   );
	FA e83(.p({r1[23][9],r1[23][10],r1[23][11]}),    .w({r1[24][11],r2[23][3]})   ); // column 23
	
	FA e84(.p({r1[24][0],r1[24][1 ],r1[24][2 ]}),    .w({r1[25][6],r2[24][0]})   );
	FA e85(.p({r1[24][3],r1[24][4 ],r1[24][5 ]}),    .w({r1[25][7],r2[24][1]})   );
	FA e86(.p({r1[24][6],r1[24][7 ],r1[24][8 ]}),    .w({r1[25][8],r2[24][2]})   );
	FA e87(.p({r1[24][9],r1[24][10],r1[24][11]}),    .w({r1[25][9],r2[24][3]})   ); // column 24
	
	assign r2[25][3] = r1[25][9];
	FA e88(.p({r1[25][0],r1[25][1],r1[25][2]}),    .w({r1[26][5],r2[25][0]})   );
	FA e89(.p({r1[25][3],r1[25][4],r1[25][5]}),    .w({r1[26][6],r2[25][1]})   );
	FA e90(.p({r1[25][6],r1[25][7],r1[25][8]}),    .w({r1[26][7],r2[25][2]})   ); // column 25

    FA e91(.p({r1[26][0],r1[26][1],r1[26][2]}),    .w({r1[27][4],r2[26][0]})   );
	FA e92(.p({r1[26][3],r1[26][4],r1[26][5]}),    .w({r1[27][5],r2[26][1]})   );
	HA e93(.p({r1[26][6],r1[26][7]}),              .w({r1[27][6],r2[26][2]})   ); // column 26
	
	assign r2[27][2] = r1[27][6];
	FA e94(.p({r1[27][0],r1[27][1],r1[27][2]}),    .w({r1[28][3],r2[27][0]})   );
	FA e95(.p({r1[27][3],r1[27][4],r1[27][5]}),    .w({r1[28][4],r2[27][1]})   ); // column 27
	
	FA e96(.p({r1[28][0],r1[28][1],r1[28][2]}),    .w({r1[29][2],r2[28][0]})   );
	HA e97(.p({r1[28][3],r1[28][4]}),              .w({r1[29][3],r2[28][1]})   ); // column 28
	
	assign r2[29][1] = r1[29][3];
	FA e98(.p({r1[29][0],r1[29][1],r1[29][2]}),    .w({r1[30][1],r2[29][0]})   ); // column 29
	
	assign r2[30][0] = r1[30][0];
	assign r2[30][1] = r1[30][1]; // column 30
	
	//////////////////////////////////////////// one more full adder stage///////////////////////
    wire r3[30:0][5:0] ; // outputs of first reduction
	wire cout;
	
	assign r3[0][0] = r2[0][0]; // column 0
	assign r3[0][1] = 1'b0; // the third reduced pp doesnt provide value
	 
	assign r3[1][0] = r2[1][0];
	assign r3[1][1] = r2[1][1]; // column 1
	
	assign r3[2][0] = r2[2][0];
	assign r3[2][1] = r2[2][1]; // column 2
	
	assign r3[3][0] = r2[3][0];
	assign r3[3][1] = r2[3][1]; // column 3
	
	assign r3[4][0] = r2[4][0];
	assign r3[4][1] = r2[4][1]; // column 4
	
	assign r3[5][0] = r2[5][0];
	assign r3[5][1] = r2[5][1]; // column 5
	
	assign r3[6][0] = r2[6][0];
	assign r3[6][1] = r2[6][1]; // column 6
	
	assign r3[7][0] = r2[7][0];
	assign r3[7][1] = r2[7][1]; // column 7
	
	assign r3[8][1] = 1'b0;
	FA e99(.p({r2[8][0],r2[8][1],r2[8][2]}),    .w({r2[9][3],r3[8][0]})   ); // column 8
	
	assign r3[9][1] = r2[9][3];
	FA e100(.p({r2[9][0],r2[9][1],r2[9][2]}),    .w({r2[10][3],r3[9][0]})   ); // column 9
	
	assign r3[10][1] = r2[10][3];
	FA e101(.p({r2[10][0],r2[10][1],r2[10][2]}),    .w({r2[11][3],r3[10][0]})   ); // column 10
	
	assign r3[11][1] = r2[11][3];
	FA e102(.p({r2[11][0],r2[11][1],r2[11][2]}),    .w({r2[12][4],r3[11][0]})   ); // column 11
	
	FA e103(.p({r2[12][0],r2[12][1],r2[12][2]}),    .w({r2[13][4],r3[12][0]})   ); 
	HA e137(.p({r2[12][3],r2[12][4]}),              .w({r2[13][5],r3[12][1]})   ); // column 12
	
	FA e104(.p({r2[13][0],r2[13][1],r2[13][2]}),    .w({r2[14][4],r3[13][0]})   );
	FA e105(.p({r2[13][3],r2[13][4],r2[13][5]}),    .w({r2[14][5],r3[13][1]})   ); // column 13
	
	FA e106(.p({r2[14][0],r2[14][1],r2[14][2]}),    .w({r2[15][4],r3[14][0]})   );
	FA e107(.p({r2[14][3],r2[14][4],r2[14][5]}),    .w({r2[15][5],r3[14][1]})   ); // column 14
	
	FA e108(.p({r2[15][0],r2[15][1],r2[15][2]}),    .w({r2[16][4],r3[15][0]})   );
	FA e109(.p({r2[15][3],r2[15][4],r2[15][5]}),    .w({r2[16][5],r3[15][1]})   ); // column 15
	
	FA e110(.p({r2[16][0],r2[16][1],r2[16][2]}),    .w({r2[17][4],r3[16][0]})   );
	FA e111(.p({r2[16][3],r2[16][4],r2[16][5]}),    .w({r2[17][5],r3[16][1]})   ); // column 16
	
	FA e112(.p({r2[17][0],r2[17][1],r2[17][2]}),    .w({r2[18][4],r3[17][0]})   );
	FA e113(.p({r2[17][3],r2[17][4],r2[17][5]}),    .w({r2[18][5],r3[17][1]})   ); // column 17
	
	FA e114(.p({r2[18][0],r2[18][1],r2[8 ][2]}),    .w({r2[19][4],r3[18][0]})   );
	FA e115(.p({r2[18][3],r2[18][4],r2[18][5]}),    .w({r2[19][5],r3[18][1]})   ); // column 18
	
	FA e116(.p({r2[19][0],r2[19][1],r2[19][2]}),    .w({r2[20][4],r3[19][0]})   );
	FA e117(.p({r2[19][3],r2[19][4],r2[19][5]}),    .w({r2[20][5],r3[19][1]})   ); // column 19
	
	FA e118(.p({r2[20][0],r2[20][1],r2[20][2]}),    .w({r2[21][4],r3[20][0]})   );
	FA e119(.p({r2[20][3],r2[20][4],r2[20][5]}),    .w({r2[21][5],r3[20][1]})   ); // column 20
	
	FA e120(.p({r2[21][0],r2[21][1],r2[21][2]}),    .w({r2[22][4],r3[21][0]})   );
	FA e121(.p({r2[21][3],r2[21][4],r2[21][5]}),    .w({r2[22][5],r3[21][1]})   ); // column 21
	
	FA e122(.p({r2[22][0],r2[22][1],r2[22][2]}),    .w({r2[23][4],r3[22][0]})   );
	FA e123(.p({r2[22][3],r2[22][4],r2[22][5]}),    .w({r2[23][5],r3[22][1]})   ); // column 22
	
	FA e124(.p({r2[23][0],r2[23][1],r2[23][2]}),    .w({r2[24][4],r3[23][0]})   );
	FA e125(.p({r2[23][3],r2[23][4],r2[23][5]}),    .w({r2[24][5],r3[23][1]})   ); // column 23
	
	FA e126(.p({r2[24][0],r2[24][1],r2[24][2]}),    .w({r2[25][4],r3[24][0]})   );
	FA e127(.p({r2[24][3],r2[24][4],r2[24][5]}),    .w({r2[25][5],r3[24][1]})   ); // column 24
	
	//assign r2[25][5] = r1[25][9];
	FA e128(.p({r2[25][0],r2[25][1],r2[25][2]}),    .w({r2[26][3],r3[25][0]})   ); 
	FA e129(.p({r2[25][3],r2[25][4],r2[25][5]}),    .w({r2[26][4],r3[25][1]})   ); // column 25
	
	FA e130(.p({r2[26][0],r2[26][1],r2[26][2]}),    .w({r2[27][3],r3[26][0]})   ); 
	HA e131(.p({r2[26][3],r2[26][4]}),              .w({r2[27][4],r3[26][1]})   ); // column 26
	
	FA e132(.p({r2[27][0],r2[27][1],r2[27][2]}),    .w({r2[28][2],r3[27][0]})   ); 
	HA e133(.p({r2[27][3],r2[27][4]}),              .w({r2[28][3],r3[27][1]})   ); // column 27
	
	assign r3[28][1] = r2[28][3];
	FA e134(.p({r2[28][0],r2[28][1],r2[28][2]}),    .w({r2[29][2],r3[28][0]})   ); // column 28
	
	assign r3[29][1] = r2[29][2];
	HA e135(.p({r2[29][0],r2[29][1]}),    .w({r2[30][2],r3[29][0]})   ); // column 29
	
	assign r3[30][1] = r2[30][2];
	HA e136(.p({r2[30][0],r2[30][1]}),    .w({cout,r3[30][0]})   ); // column 30
//	assign r3[29][1] = 1'b0;
//	FA e135(.p({r2[29][0],r2[29][1],r2[29][2]}),    .w({r2[30][2],r3[29][0]})   ); // column 29
	
//	assign r3[30][1] = 1'b0;
//	FA e136(.p({r2[30][0],r2[30][1],r2[30][2]}),    .w({cout,r3[30][0]})   ); // column 30
	
	//////////////////////////////////////////// Outputs of processing block   ////////////////////////
	assign out1[0] = r3[0][0];    
    assign out1[1] = r3[1][0];
    assign out1[2] = r3[2][0];
    assign out1[3] = r3[3][0];
    assign out1[4] = r3[4][0];
    assign out1[5] = r3[5][0];
    assign out1[6] = r3[6][0];
    assign out1[7] = r3[7][0];
    assign out1[8] = r3[8][0];
    assign out1[9] = r3[9][0];
    assign out1[10] = r3[10][0];
    assign out1[11] = r3[11][0];
    assign out1[12] = r3[12][0];
    assign out1[13] = r3[13][0];
    assign out1[14] = r3[14][0];
	assign out1[15] = r3[15][0];
    assign out1[16] = r3[16][0];
    assign out1[17] = r3[17][0];
    assign out1[18] = r3[18][0];
    assign out1[19] = r3[19][0];
	assign out1[20] = r3[20][0];
	assign out1[21] = r3[21][0];
    assign out1[22] = r3[22][0];
    assign out1[23] = r3[23][0];
    assign out1[24] = r3[24][0];
    assign out1[25] = r3[25][0];
    assign out1[26] = r3[26][0];
    assign out1[27] = r3[27][0];
    assign out1[28] = r3[28][0];
    assign out1[29] = r3[29][0];
    assign out1[30] = r3[30][0];
    
    assign out2[0] = r3[0][1];    
    assign out2[1] = r3[1][1];
    assign out2[2] = r3[2][1];
    assign out2[3] = r3[3][1];
    assign out2[4] = r3[4][1];
    assign out2[5] = r3[5][1];
    assign out2[6] = r3[6][1];
    assign out2[7] = r3[7][1];
    assign out2[8] = r3[8][1];
    assign out2[9] = r3[9][1];
    assign out2[10] = r3[10][1];
    assign out2[11] = r3[11][1];
    assign out2[12] = r3[12][1];
    assign out2[13] = r3[13][1];
    assign out2[14] = r3[14][1];
	assign out2[15] = r3[15][1];
    assign out2[16] = r3[16][1];
    assign out2[17] = r3[17][1];
    assign out2[18] = r3[18][1];
    assign out2[19] = r3[19][1];
	assign out2[20] = r3[20][1];
	assign out2[21] = r3[21][1];
    assign out2[22] = r3[22][1];
    assign out2[23] = r3[23][1];
    assign out2[24] = r3[24][1];
    assign out2[25] = r3[25][1];
    assign out2[26] = r3[26][1];
    assign out2[27] = r3[27][1];
    assign out2[28] = r3[28][1];
    assign out2[29] = r3[29][1];
    assign out2[30] = r3[30][1];

endmodule

////////////////////////////////////////////// 16 bit 2 step processing block //////////////////////
module processing_block_16_2step(
input p[15:0][15:0],
output [30:0]out1,
output [30:0]out2);
      
    ////////////////////////////////////////// PP REDUCTION STEP ONE   ////////////////////////  
    wire r1[30:0][7:0] ; // outputs of first reduction
    
    assign r1[0][0] = p[0][0];                                                 // column 0
    assign r1[1][0] = p[1][0]; assign r1[1][1] = p[0][1];                       // column 1
    compressor3_2 c1   (.p({p[2][0]  ,p[1][1]  ,p[0][2]}),                                                                                                                    .w({r1[2][0] ,r1[2][1]}));                                                // column 2
    compressor4_2 c2   (.p({p[3][0]  ,p[2][1]  ,p[1][2] ,p[0][3]}),                                                                                                           .w({r1[3][0] ,r1[3][1]}));                                              // column 3
    compressor5_3 c3   (.p({p[4][0]  ,p[3][1]  ,p[2][2] ,p[1][3] ,p[0][4]}),                                                                                                  .w({r1[4][0] ,r1[4][1] ,r1[4][2]}));                                      // column 4
    compressor6_3 c4   (.p({p[5][0]  ,p[4][1]  ,p[3][2] ,p[2][3] ,p[1][4]  ,p[0][5]}),                                                                                        .w({r1[5][0] ,r1[5][1] ,r1[5][2]}));                                    // column 5
    compressor7_4 c5   (.p({p[6][0]  ,p[5][1]  ,p[4][2] ,p[3][3] ,p[2][4]  ,p[1][5] ,p[0][6]}),                                                                               .w({r1[6][0] ,r1[6][1] ,r1[6][2] ,r1[6][3]}));                               // column 6
    compressor8_4 c6   (.p({p[7][0]  ,p[6][1]  ,p[5][2] ,p[4][3] ,p[3][4]  ,p[2][5] ,p[1][6],p[0][7]}),                                                                       .w({r1[7][0] ,r1[7][1] ,r1[7][2] ,r1[7][3]}));                                // column 7
    compressor9_5 c7   (.p({p[8][0]  ,p[7][1]  ,p[6][2] ,p[5][3] ,p[4][4]  ,p[3][5] ,p[2][6],p[1][7],p[0][8]}),                                                               .w({r1[8][0] ,r1[8][1] ,r1[8][2] ,r1[8][3] ,r1[8][4]}));                       // column 8
    compressor10_5 c8  (.p({p[9][0]  ,p[8][1]  ,p[7][2] ,p[6][3] ,p[5][4]  ,p[4][5] ,p[3][6],p[2][7],p[1][8],p[0][9]}),                                                       .w({r1[9][0] ,r1[9][1] ,r1[9][2] ,r1[9][3] ,r1[9][4]}));                         // column 9
    compressor11_6 c9  (.p({p[10][0] ,p[9][1]  ,p[8][2] ,p[7][3] ,p[6][4]  ,p[5][5] ,p[4][6],p[3][7],p[2][8],p[1][9],p[0][10]}),                                              .w({r1[10][0],r1[10][1],r1[10][2],r1[10][3],r1[10][4],r1[10][5]}));              // column 10
    compressor12_6 c10 (.p({p[11][0] ,p[10][1] ,p[9][2] ,p[8][3] ,p[7][4]  ,p[6][5] ,p[5][6],p[4][7],p[3][8],p[2][9],p[1][10],p[0][11]}),                                     .w({r1[11][0],r1[11][1],r1[11][2],r1[11][3],r1[11][4],r1[11][5]}));              // column 11
    compressor13_7 c11 (.p({p[12][0] ,p[11][1] ,p[10][2],p[9][3] ,p[8][4]  ,p[7][5] ,p[6][6],p[5][7],p[4][8],p[3][9],p[2][10],p[1][11],p[0][12]}),                            .w({r1[12][0],r1[12][1],r1[12][2],r1[12][3],r1[12][4],r1[12][5],r1[12][6]}));     // column 12
    compressor14_7 c12 (.p({p[13][0] ,p[12][1] ,p[11][2],p[10][3],p[9][4]  ,p[8][5] ,p[7][6],p[6][7],p[5][8],p[4][9],p[3][10],p[2][11],p[1][12],p[0][13]}),                   .w({r1[13][0],r1[13][1],r1[13][2],r1[13][3],r1[13][4],r1[13][5],r1[13][6]}));      // column 13
    compressor15_8 c13 (.p({p[14][0] ,p[13][1] ,p[12][2],p[11][3],p[10][4] ,p[9][5] ,p[8][6],p[7][7],p[6][8],p[5][9],p[4][10],p[3][11],p[2][12],p[1][13],p[0][14]}),          .w({r1[14][0],r1[14][1],r1[14][2],r1[14][3],r1[14][4],r1[14][5],r1[14][6],r1[14][7]})); // column 14
    compressor16_8 c14 (.p({p[15][0] ,p[14][1] ,p[13][2],p[12][3],p[11][4] ,p[10][5],p[9][6],p[8][7],p[7][8],p[6][9],p[5][10],p[4][11],p[3][12],p[2][13],p[1][14],p[0][15]}), .w({r1[15][0],r1[15][1],r1[15][2],r1[15][3],r1[15][4],r1[15][5],r1[15][6],r1[15][7]})); // column 15
    
    compressor14_7 c15 (.p({p[15][1] ,p[14][2] ,p[13][3],p[12][4],p[11][5]  ,p[10][6] ,p[9][7],p[8][8],p[7][9],p[6][10],p[5][11],p[4][12],p[3][13],p[2][14]}),                .w({r1[16][0],r1[16][1],r1[16][2],r1[16][3],r1[16][4],r1[16][5],r1[16][6]}));
    assign r1[16][7] = p[1][15];// column 16
    
    FA e1(.p({p[15][2],p[14][3],p[13][4]}), .w({r1[18][0],r1[17][0]})   );
    FA e2(.p({p[12][5],p[11][6],p[10][7]}), .w({r1[18][1],r1[17][1]})   );
    FA e3(.p({p[9][8],p[8][9],p[7][10]}), .w({r1[18][2],r1[17][2]})   ); 
    assign r1[17][3] = p[6][11];
    assign r1[17][4] = p[5][12];
    assign r1[17][5] = p[4][13];
    assign r1[17][6] = p[3][14];
    assign r1[17][7] = p[2][15];//column 17
    
    FA e4(.p({p[15][3],p[14][4],p[13][5]}), .w({r1[19][0],r1[18][3]})   );
    FA e5(.p({p[12][6],p[11][7],p[10][8]}), .w({r1[19][1],r1[18][4]})   );
    FA e6(.p({p[9][9],p[8][10],p[7][11]}), .w({r1[19][2],r1[18][5]})   ); 
    FA e7(.p({p[6][12],p[5][13],p[4][14]}), .w({r1[19][3],r1[18][6]})   );
    assign r1[18][7] = p[3][15]; //column 18
    
    FA e8(.p({p[15][4],p[14][5],p[13][6]}),  .w({r1[20][0],r1[19][4]})   );
    FA e9(.p({p[12][7],p[11][8],p[10][9]}),  .w({r1[20][1],r1[19][5]})   );
    FA e10(.p({p[9][10],p[8][11],p[7][12]}), .w({r1[20][2],r1[19][6]})   ); 
    FA e11(.p({p[6][13],p[5][14],p[4][15]}), .w({r1[20][3],r1[19][7]})   ); //column 19
    
    FA e12(.p({p[15][5],p[14][6],p[13][7]}),  .w({r1[21][0],r1[20][4]})   );
    FA e13(.p({p[12][8],p[11][9],p[10][10]}), .w({r1[21][1],r1[20][5]})   );
    FA e14(.p({p[9][11],p[8][12],p[7][13]}),  .w({r1[21][2],r1[20][6]})   );
    HA e15(.p({p[6][14],p[5][15]}),           .w({r1[21][3],r1[20][7]})   ); //column 20
    
    FA e16(.p({p[15][6],p[14][7],p[13][8]}),   .w({r1[22][0],r1[21][4]})   );
    FA e17(.p({p[12][9],p[11][10],p[10][11]}), .w({r1[22][1],r1[21][5]})   );
    FA e18(.p({p[9][12],p[8][13],p[7][14]}),   .w({r1[22][2],r1[21][6]})   );
    assign r1[21][7] = p[6][15]; //column 21
    
    FA e19(.p({p[15][7],p[14][8],p[13][9]}),    .w({r1[23][0],r1[22][3]})   );
    FA e20(.p({p[12][10],p[11][11],p[10][12]}), .w({r1[23][1],r1[22][4]})   ); 
    assign r1[22][5] = p[9][13];
    assign r1[22][6] = p[8][14];
    assign r1[22][7] = p[7][15]; //column 22
    
    FA e21(.p({p[15][8],p[14][9],p[13][10]}), .w({r1[24][0],r1[23][2]})   );
    assign r1[23][3] = p[12][11];
    assign r1[23][4] = p[11][12];
    assign r1[23][5] = p[10][13];
    assign r1[23][6] = p[9][14];
    assign r1[23][7] = p[8][15]; //column 23
    
    assign r1[24][1] = p[15][9];
    assign r1[24][2] = p[14][10];
    assign r1[24][3] = p[13][11];
    assign r1[24][4] = p[12][12];
    assign r1[24][5] = p[11][13];
    assign r1[24][6] = p[10][14];
    assign r1[24][7] = p[9][15]; //column 24
    
    assign r1[25][0] = p[15][10];
    assign r1[25][1] = p[14][11];
    assign r1[25][2] = p[13][12];
    assign r1[25][3] = p[12][13];
    assign r1[25][4] = p[11][14];
    assign r1[25][5] = p[10][15]; //column 25
    
    assign r1[26][0] = p[15][11];
    assign r1[26][1] = p[14][12];
    assign r1[26][2] = p[13][13];
    assign r1[26][3] = p[12][14];
    assign r1[26][4] = p[11][15]; //column 26
    
    assign r1[27][0] = p[15][12];
    assign r1[27][1] = p[14][13];
    assign r1[27][2] = p[13][14];
    assign r1[27][3] = p[12][15]; //column 27
    
    assign r1[28][0] = p[15][13];
    assign r1[28][1] = p[14][14];
    assign r1[28][2] = p[13][15]; //column 28
    
    assign r1[29][0] = p[15][14];
    assign r1[29][1] = p[14][15]; //column 29
   
    assign r1[30][0] = p[15][15]; //column 30
    
    
    ////////////////////////////////////////// PP REDUCTION STEP TWO   ////////////////////////  
    wire r2[30:0][5:0] ; // outputs of first reduction
    
    assign r2[0][0] = r1[0][0];// column 0
    
    assign r2[1][0] = r1[1][0];
    assign r2[1][1] = r1[1][1];// column 1
    
    assign r2[2][0] = r1[2][0];
    assign r2[2][1] = r1[2][1];// column 2
    
    assign r2[3][0] = r1[3][0];
    assign r2[3][1] = r1[3][1];// column 3
    
    compressor3_2 c16   (.p({r1[4][0]   ,r1[4][1]   ,r1[4][2]}),                                                       .w({r2[4][0]  ,r2[4][1]})); // column 4
    compressor3_2 c17   (.p({r1[5][0]   ,r1[5][1]   ,r1[5][2]}),                                                       .w({r2[5][0]  ,r2[5][1]})); // column 5
    compressor4_2 c18   (.p({r1[6][0]   ,r1[6][1]   ,r1[6][2]  ,r1[6][3]}),                                            .w({r2[6][0]  ,r2[6][1]})); // column 6
    compressor4_2 c19   (.p({r1[7][0]   ,r1[7][1]   ,r1[7][2]  ,r1[7][3]}),                                            .w({r2[7][0]  ,r2[7][1]})); // column 7
    compressor5_3 c20   (.p({r1[8][0]   ,r1[8][1]   ,r1[8][2]  ,r1[8][3]  ,r1[8][4]}),                                 .w({r2[8][0]  ,r2[8][1] ,r2[8][2]})); // column 8
    compressor5_3 c21   (.p({r1[9][0]   ,r1[9][1]   ,r1[9][2]  ,r1[9][3]  ,r1[9][4]}),                                 .w({r2[9][0]  ,r2[9][1] ,r2[9][2]})); // column 9
    compressor6_3 c22   (.p({r1[10][0]  ,r1[10][1]  ,r1[10][2] ,r1[10][3] ,r1[10][4],r1[10][5]}),                      .w({r2[10][0] ,r2[10][1],r2[10][2]})); // column 10
    compressor6_3 c23   (.p({r1[11][0]  ,r1[11][1]  ,r1[11][2] ,r1[11][3] ,r1[11][4],r1[11][5]}),                      .w({r2[11][0] ,r2[11][1],r2[11][2]})); // column 11
    compressor7_4 c24   (.p({r1[12][0]  ,r1[12][1]  ,r1[12][2] ,r1[12][3] ,r1[12][4],r1[12][5],r1[12][6]}),            .w({r2[12][0] ,r2[12][1],r2[12][2],r2[12][3]})); // column 12
    compressor7_4 c25   (.p({r1[13][0]  ,r1[13][1]  ,r1[13][2] ,r1[13][3] ,r1[13][4],r1[13][5],r1[13][6]}),            .w({r2[13][0] ,r2[13][1],r2[13][2],r2[13][3]})); // column 13
    compressor8_4 c26   (.p({r1[14][0]  ,r1[14][1]  ,r1[14][2] ,r1[14][3] ,r1[14][4],r1[14][5],r1[14][6],r1[14][7]}),  .w({r2[14][0] ,r2[14][1],r2[14][2],r2[14][3]})); // column 14
    compressor8_4 c27   (.p({r1[15][0]  ,r1[15][1]  ,r1[15][2] ,r1[15][3] ,r1[15][4],r1[15][5],r1[15][6],r1[15][7]}),  .w({r2[15][0] ,r2[15][1],r2[15][2],r2[15][3]})); // column 15
    compressor8_4 c28   (.p({r1[16][0]  ,r1[16][1]  ,r1[16][2] ,r1[16][3] ,r1[16][4],r1[16][5],r1[16][6],r1[16][7]}),  .w({r2[16][0] ,r2[16][1],r2[16][2],r2[16][3]})); // column 16
    compressor8_4 c29   (.p({r1[17][0]  ,r1[17][1]  ,r1[17][2] ,r1[17][3] ,r1[17][4],r1[17][5],r1[17][6],r1[17][7]}),  .w({r2[17][0] ,r2[17][1],r2[17][2],r2[17][3]})); // column 17
    compressor8_4 c30   (.p({r1[18][0]  ,r1[18][1]  ,r1[18][2] ,r1[18][3] ,r1[18][4],r1[18][5],r1[18][6],r1[18][7]}),  .w({r2[18][0] ,r2[18][1],r2[18][2],r2[18][3]})); // column 18
    compressor8_4 c31   (.p({r1[19][0]  ,r1[19][1]  ,r1[19][2] ,r1[19][3] ,r1[19][4],r1[19][5],r1[19][6],r1[19][7]}),  .w({r2[19][0] ,r2[19][1],r2[19][2],r2[19][3]})); // column 19
    compressor8_4 c32   (.p({r1[20][0]  ,r1[20][1]  ,r1[20][2] ,r1[20][3] ,r1[20][4],r1[20][5],r1[20][6],r1[20][7]}),  .w({r2[20][0] ,r2[20][1],r2[20][2],r2[20][3]})); // column 20
    compressor8_4 c33   (.p({r1[21][0]  ,r1[21][1]  ,r1[21][2] ,r1[21][3] ,r1[21][4],r1[21][5],r1[21][6],r1[21][7]}),  .w({r2[21][0] ,r2[21][1],r2[21][2],r2[21][3]})); // column 21
    compressor8_4 c34   (.p({r1[22][0]  ,r1[22][1]  ,r1[22][2] ,r1[22][3] ,r1[22][4],r1[22][5],r1[22][6],r1[22][7]}),  .w({r2[22][0] ,r2[22][1],r2[22][2],r2[22][3]})); // column 22
    compressor8_4 c35   (.p({r1[23][0]  ,r1[23][1]  ,r1[23][2] ,r1[23][3] ,r1[23][4],r1[23][5],r1[23][6],r1[23][7]}),  .w({r2[23][0] ,r2[23][1],r2[23][2],r2[23][3]})); // column 23
    
    FA e22(.p({r1[24][0],r1[24][1],r1[24][2]}), .w({r2[25][0],r2[24][0]})   );
    FA e23(.p({r1[24][3],r1[24][4],r1[24][5]}), .w({r2[25][1],r2[24][1]})   ); 
    assign r2[24][2] = r1[24][6];
    assign r2[24][3] = r1[24][7]; // column 24
    
    FA e24(.p({r1[25][0],r1[25][1],r1[25][2]}), .w({r2[26][0],r2[25][2]})   );
    FA e25(.p({r1[25][3],r1[25][4],r1[25][5]}), .w({r2[26][1],r2[25][3]})   ); // column 25
    
    FA e26(.p({r1[26][0],r1[26][1],r1[26][2]}), .w({r2[27][0],r2[26][2]})   );
    HA e27(.p({r1[26][3],r1[26][4]}),           .w({r2[27][1],r2[26][3]})   ); // column 26
    
    FA e28(.p({r1[27][0],r1[27][1],r1[27][2]}), .w({r2[28][0],r2[27][2]})   ); 
    assign r2[27][3] = r1[27][3]; // column 27
						
    assign r2[28][1] = r1[28][0];
    assign r2[28][2] = r1[28][1];
    assign r2[28][3] = r1[28][2]; //column 28
						
    assign r2[29][0] = r1[29][0];
    assign r2[29][1] = r1[29][1]; //column 29
						
    assign r2[30][0] = r1[30][0]; //column 30
    
    ////////////////////////////////////////////////////// Exact adders //////////////////////////////////////////
    wire r3[30:0][1:0] ;
    
    assign r3[0][0] = r2[0][0];// column 0
    assign r3[0][1] = 1'b0; // the third reduced pp doesnt provide value
    
    assign r3[1][0] = r2[1][0];
    assign r3[1][1] = r2[1][1];// column 1
    
    assign r3[2][0] = r2[2][0];
    assign r3[2][1] = r2[2][1];// column 2
    
    assign r3[3][0] = r2[3][0];
    assign r3[3][1] = r2[3][1];// column 3
    
    assign r3[4][0] = r2[4][0];
    assign r3[4][1] = r2[4][1];// column 4
    
    assign r3[5][0] = r2[5][0];
    assign r3[5][1] = r2[5][1];// column 5
    
    assign r3[6][0] = r2[6][0];
    assign r3[6][1] = r2[6][1];// column 6
	
	assign r3[7][0] = r2[7][0];
    assign r3[7][1] = r2[7][1];// column 7
    
    assign r3[8][1] = 1'b0;
    FA e29(.p({r2[8][0],r2[8][1],r2[8][2]}), .w({r2[9][3],r3[8][0]})   ); // column 8
    
    assign r3[9][1] = r2[9][3];
    FA e30(.p({r2[9][0],r2[9][1],r2[9][2]}), .w({r2[10][3],r3[9][0]})   ); // column 9
    
    assign r3[10][1] = r2[10][3];
    FA e31(.p({r2[10][0],r2[10][1],r2[10][2]}), .w({r2[11][3],r3[10][0]})   ); // column 10
    
    assign r3[11][1] = r2[11][3];
    FA e32(.p({r2[11][0],r2[11][1],r2[11][2]}), .w({r2[12][4],r3[11][0]})   ); // column 11
    
    HA e33(.p({r2[12][3],r2[12][4]}), .w({r2[13][5],r3[12][1]})   ); 
    FA e34(.p({r2[12][0],r2[12][1],r2[12][2]}), .w({r2[13][4],r3[12][0]})   ); // column 12
    
    FA e35(.p({r2[13][0],r2[13][1],r2[13][2]}), .w({r2[14][4],r3[13][0]})   ); 
    FA e36(.p({r2[13][3],r2[13][4],r2[13][5]}), .w({r2[14][5],r3[13][1]})   ); // column 13
    FA e37(.p({r2[14][0],r2[14][1],r2[14][2]}), .w({r2[15][4],r3[14][0]})   ); 
    FA e38(.p({r2[14][3],r2[14][4],r2[14][5]}), .w({r2[15][5],r3[14][1]})   ); // column 14
    FA e39(.p({r2[15][0],r2[15][1],r2[15][2]}), .w({r2[16][4],r3[15][0]})   ); 
    FA e40(.p({r2[15][3],r2[15][4],r2[15][5]}), .w({r2[16][5],r3[15][1]})   ); // column 15
    FA e41(.p({r2[16][0],r2[16][1],r2[16][2]}), .w({r2[17][4],r3[16][0]})   ); 
    FA e42(.p({r2[16][3],r2[16][4],r2[16][5]}), .w({r2[17][5],r3[16][1]})   ); // column 16
    FA e43(.p({r2[17][0],r2[17][1],r2[17][2]}), .w({r2[18][4],r3[17][0]})   ); 
    FA e44(.p({r2[17][3],r2[17][4],r2[17][5]}), .w({r2[18][5],r3[17][1]})   ); // column 17
    FA e45(.p({r2[18][0],r2[18][1],r2[18][2]}), .w({r2[19][4],r3[18][0]})   ); 
    FA e46(.p({r2[18][3],r2[18][4],r2[18][5]}), .w({r2[19][5],r3[18][1]})   ); // column 18
    FA e47(.p({r2[19][0],r2[19][1],r2[19][2]}), .w({r2[20][4],r3[19][0]})   ); 
    FA e48(.p({r2[19][3],r2[19][4],r2[19][5]}), .w({r2[20][5],r3[19][1]})   ); // column 19
    FA e49(.p({r2[20][0],r2[20][1],r2[20][2]}), .w({r2[21][4],r3[20][0]})   ); 
    FA e50(.p({r2[20][3],r2[20][4],r2[20][5]}), .w({r2[21][5],r3[20][1]})   ); // column 20
    FA e51(.p({r2[21][0],r2[21][1],r2[21][2]}), .w({r2[22][4],r3[21][0]})   ); 
    FA e52(.p({r2[21][3],r2[21][4],r2[21][5]}), .w({r2[22][5],r3[21][1]})   ); // column 21
    FA e53(.p({r2[22][0],r2[22][1],r2[22][2]}), .w({r2[23][4],r3[22][0]})   ); 
    FA e54(.p({r2[22][3],r2[22][4],r2[22][5]}), .w({r2[23][5],r3[22][1]})   ); // column 22
    FA e55(.p({r2[23][0],r2[23][1],r2[23][2]}), .w({r2[24][4],r3[23][0]})   ); 
    FA e56(.p({r2[23][3],r2[23][4],r2[23][5]}), .w({r2[24][5],r3[23][1]})   ); // column 23
    FA e57(.p({r2[24][0],r2[24][1],r2[24][2]}), .w({r2[25][4],r3[24][0]})   ); 
    FA e58(.p({r2[24][3],r2[24][4],r2[24][5]}), .w({r2[25][5],r3[24][1]})   ); // column 24
    FA e59(.p({r2[25][0],r2[25][1],r2[25][2]}), .w({r2[26][4],r3[25][0]})   ); 
    FA e60(.p({r2[25][3],r2[25][4],r2[25][5]}), .w({r2[26][5],r3[25][1]})   ); // column 25
    FA e61(.p({r2[26][0],r2[26][1],r2[26][2]}), .w({r2[27][4],r3[26][0]})   ); 
    FA e62(.p({r2[26][3],r2[26][4],r2[26][5]}), .w({r2[27][5],r3[26][1]})   ); // column 26
    FA e63(.p({r2[27][0],r2[27][1],r2[27][2]}), .w({r2[28][4],r3[27][0]})   ); 
    FA e64(.p({r2[27][3],r2[27][4],r2[27][5]}), .w({r2[28][5],r3[27][1]})   ); // column 27
    FA e65(.p({r2[28][0],r2[28][1],r2[28][2]}), .w({r2[29][2],r3[28][0]})   ); 
    FA e66(.p({r2[28][3],r2[28][4],r2[28][5]}), .w({r2[29][3],r3[28][1]})   ); // column 28
    
    assign r3[29][1] = r2[29][3];
    FA e67(.p({r2[29][0],r2[29][1],r2[29][2]}), .w({r2[30][1],r3[29][0]})   ); // column 29
    
    assign r3[30][0] = r2[30][0];
    assign r3[30][1] = r2[30][1]; // column 30

    //////////////////////////////////////////// Outputs of processing block   ////////////////////////
	assign out1[0] = r3[0][0];    
    assign out1[1] = r3[1][0];
    assign out1[2] = r3[2][0];
    assign out1[3] = r3[3][0];
    assign out1[4] = r3[4][0];
    assign out1[5] = r3[5][0];
    assign out1[6] = r3[6][0];
    assign out1[7] = r3[7][0];
    assign out1[8] = r3[8][0];
    assign out1[9] = r3[9][0];
    assign out1[10] = r3[10][0];
    assign out1[11] = r3[11][0];
    assign out1[12] = r3[12][0];
    assign out1[13] = r3[13][0];
    assign out1[14] = r3[14][0];
	assign out1[15] = r3[15][0];
    assign out1[16] = r3[16][0];
    assign out1[17] = r3[17][0];
    assign out1[18] = r3[18][0];
    assign out1[19] = r3[19][0];
	assign out1[20] = r3[20][0];
	assign out1[21] = r3[21][0];
    assign out1[22] = r3[22][0];
    assign out1[23] = r3[23][0];
    assign out1[24] = r3[24][0];
    assign out1[25] = r3[25][0];
    assign out1[26] = r3[26][0];
    assign out1[27] = r3[27][0];
    assign out1[28] = r3[28][0];
    assign out1[29] = r3[29][0];
    assign out1[30] = r3[30][0];
    
    assign out2[0] = r3[0][1];    
    assign out2[1] = r3[1][1];
    assign out2[2] = r3[2][1];
    assign out2[3] = r3[3][1];
    assign out2[4] = r3[4][1];
    assign out2[5] = r3[5][1];
    assign out2[6] = r3[6][1];
    assign out2[7] = r3[7][1];
    assign out2[8] = r3[8][1];
    assign out2[9] = r3[9][1];
    assign out2[10] = r3[10][1];
    assign out2[11] = r3[11][1];
    assign out2[12] = r3[12][1];
    assign out2[13] = r3[13][1];
    assign out2[14] = r3[14][1];
	assign out2[15] = r3[15][1];
    assign out2[16] = r3[16][1];
    assign out2[17] = r3[17][1];
    assign out2[18] = r3[18][1];
    assign out2[19] = r3[19][1];
	assign out2[20] = r3[20][1];
	assign out2[21] = r3[21][1];
    assign out2[22] = r3[22][1];
    assign out2[23] = r3[23][1];
    assign out2[24] = r3[24][1];
    assign out2[25] = r3[25][1];
    assign out2[26] = r3[26][1];
    assign out2[27] = r3[27][1];
    assign out2[28] = r3[28][1];
    assign out2[29] = r3[29][1];
    assign out2[30] = r3[30][1];

 endmodule
 
 
////////////////////////////////////////////// 16 bit 3 step processing block //////////////////////
module processing_block_16_3step(
input p[15:0][15:0],
output [30:0]out1,
output [30:0]out2
    );  

    ////////////////////////////////////////// PP REDUCTION STEP ONE   ////////////////////////  
    wire r1[30:0][7:0] ; // outputs of first reduction
    
    assign r1[0][0] = p[0][0];                                                 // column 0
    assign r1[1][0] = p[1][0]; assign r1[1][1] = p[0][1];                       // column 1
    compressor3_2 c1   (.p({p[2][0]  ,p[1][1]  ,p[0][2]}),                                                                                                                    .w({r1[2][0] ,r1[2][1]}));                                                // column 2
    compressor4_2 c2   (.p({p[3][0]  ,p[2][1]  ,p[1][2] ,p[0][3]}),                                                                                                           .w({r1[3][0] ,r1[3][1]}));                                              // column 3
    compressor5_3 c3   (.p({p[4][0]  ,p[3][1]  ,p[2][2] ,p[1][3] ,p[0][4]}),                                                                                                  .w({r1[4][0] ,r1[4][1] ,r1[4][2]}));                                      // column 4
    compressor6_3 c4   (.p({p[5][0]  ,p[4][1]  ,p[3][2] ,p[2][3] ,p[1][4]  ,p[0][5]}),                                                                                        .w({r1[5][0] ,r1[5][1] ,r1[5][2]}));                                    // column 5
    compressor7_4 c5   (.p({p[6][0]  ,p[5][1]  ,p[4][2] ,p[3][3] ,p[2][4]  ,p[1][5] ,p[0][6]}),                                                                               .w({r1[6][0] ,r1[6][1] ,r1[6][2] ,r1[6][3]}));                               // column 6
    compressor8_4 c6   (.p({p[7][0]  ,p[6][1]  ,p[5][2] ,p[4][3] ,p[3][4]  ,p[2][5] ,p[1][6],p[0][7]}),                                                                       .w({r1[7][0] ,r1[7][1] ,r1[7][2] ,r1[7][3]}));                                // column 7
    compressor9_5 c7   (.p({p[8][0]  ,p[7][1]  ,p[6][2] ,p[5][3] ,p[4][4]  ,p[3][5] ,p[2][6],p[1][7],p[0][8]}),                                                               .w({r1[8][0] ,r1[8][1] ,r1[8][2] ,r1[8][3] ,r1[8][4]}));                       // column 8
    compressor10_5 c8  (.p({p[9][0]  ,p[8][1]  ,p[7][2] ,p[6][3] ,p[5][4]  ,p[4][5] ,p[3][6],p[2][7],p[1][8],p[0][9]}),                                                       .w({r1[9][0] ,r1[9][1] ,r1[9][2] ,r1[9][3] ,r1[9][4]}));                         // column 9
    compressor11_6 c9  (.p({p[10][0] ,p[9][1]  ,p[8][2] ,p[7][3] ,p[6][4]  ,p[5][5] ,p[4][6],p[3][7],p[2][8],p[1][9],p[0][10]}),                                              .w({r1[10][0],r1[10][1],r1[10][2],r1[10][3],r1[10][4],r1[10][5]}));              // column 10
    compressor12_6 c10 (.p({p[11][0] ,p[10][1] ,p[9][2] ,p[8][3] ,p[7][4]  ,p[6][5] ,p[5][6],p[4][7],p[3][8],p[2][9],p[1][10],p[0][11]}),                                     .w({r1[11][0],r1[11][1],r1[11][2],r1[11][3],r1[11][4],r1[11][5]}));              // column 11
    compressor13_7 c11 (.p({p[12][0] ,p[11][1] ,p[10][2],p[9][3] ,p[8][4]  ,p[7][5] ,p[6][6],p[5][7],p[4][8],p[3][9],p[2][10],p[1][11],p[0][12]}),                            .w({r1[12][0],r1[12][1],r1[12][2],r1[12][3],r1[12][4],r1[12][5],r1[12][6]}));     // column 12
    compressor14_7 c12 (.p({p[13][0] ,p[12][1] ,p[11][2],p[10][3],p[9][4]  ,p[8][5] ,p[7][6],p[6][7],p[5][8],p[4][9],p[3][10],p[2][11],p[1][12],p[0][13]}),                   .w({r1[13][0],r1[13][1],r1[13][2],r1[13][3],r1[13][4],r1[13][5],r1[13][6]}));      // column 13
    compressor15_8 c13 (.p({p[14][0] ,p[13][1] ,p[12][2],p[11][3],p[10][4] ,p[9][5] ,p[8][6],p[7][7],p[6][8],p[5][9],p[4][10],p[3][11],p[2][12],p[1][13],p[0][14]}),          .w({r1[14][0],r1[14][1],r1[14][2],r1[14][3],r1[14][4],r1[14][5],r1[14][6],r1[14][7]})); // column 14
    compressor16_8 c14 (.p({p[15][0] ,p[14][1] ,p[13][2],p[12][3],p[11][4] ,p[10][5],p[9][6],p[8][7],p[7][8],p[6][9],p[5][10],p[4][11],p[3][12],p[2][13],p[1][14],p[0][15]}), .w({r1[15][0],r1[15][1],r1[15][2],r1[15][3],r1[15][4],r1[15][5],r1[15][6],r1[15][7]})); // column 15
    
    compressor14_7 c15 (.p({p[15][1] ,p[14][2] ,p[13][3],p[12][4],p[11][5]  ,p[10][6] ,p[9][7],p[8][8],p[7][9],p[6][10],p[5][11],p[4][12],p[3][13],p[2][14]}),                .w({r1[16][0],r1[16][1],r1[16][2],r1[16][3],r1[16][4],r1[16][5],r1[16][6]}));
    assign r1[16][7] = p[1][15];// column 16
    
    FA e1(.p({p[15][2],p[14][3],p[13][4]}), .w({r1[18][0],r1[17][0]})   );
    FA e2(.p({p[12][5],p[11][6],p[10][7]}), .w({r1[18][1],r1[17][1]})   );
    FA e3(.p({p[9][8],p[8][9],p[7][10]}), .w({r1[18][2],r1[17][2]})   ); 
    assign r1[17][3] = p[6][11];
    assign r1[17][4] = p[5][12];
    assign r1[17][5] = p[4][13];
    assign r1[17][6] = p[3][14];
    assign r1[17][7] = p[2][15];//column 17
    
    FA e4(.p({p[15][3],p[14][4],p[13][5]}), .w({r1[19][0],r1[18][3]})   );
    FA e5(.p({p[12][6],p[11][7],p[10][8]}), .w({r1[19][1],r1[18][4]})   );
    FA e6(.p({p[9][9],p[8][10],p[7][11]}), .w({r1[19][2],r1[18][5]})   ); 
    FA e7(.p({p[6][12],p[5][13],p[4][14]}), .w({r1[19][3],r1[18][6]})   );
    assign r1[18][7] = p[3][15]; //column 18
    
    FA e8(.p({p[15][4],p[14][5],p[13][6]}),  .w({r1[20][0],r1[19][4]})   );
    FA e9(.p({p[12][7],p[11][8],p[10][9]}),  .w({r1[20][1],r1[19][5]})   );
    FA e10(.p({p[9][10],p[8][11],p[7][12]}), .w({r1[20][2],r1[19][6]})   ); 
    FA e11(.p({p[6][13],p[5][14],p[4][15]}), .w({r1[20][3],r1[19][7]})   ); //column 19
    
    FA e12(.p({p[15][5],p[14][6],p[13][7]}),  .w({r1[21][0],r1[20][4]})   );
    FA e13(.p({p[12][8],p[11][9],p[10][10]}), .w({r1[21][1],r1[20][5]})   );
    FA e14(.p({p[9][11],p[8][12],p[7][13]}),  .w({r1[21][2],r1[20][6]})   );
    HA e15(.p({p[6][14],p[5][15]}),           .w({r1[21][3],r1[20][7]})   ); //column 20
    
    FA e16(.p({p[15][6],p[14][7],p[13][8]}),   .w({r1[22][0],r1[21][4]})   );
    FA e17(.p({p[12][9],p[11][10],p[10][11]}), .w({r1[22][1],r1[21][5]})   );
    FA e18(.p({p[9][12],p[8][13],p[7][14]}),   .w({r1[22][2],r1[21][6]})   );
    assign r1[21][7] = p[6][15]; //column 21
    
    FA e19(.p({p[15][7],p[14][8],p[13][9]}),    .w({r1[23][0],r1[22][3]})   );
    FA e20(.p({p[12][10],p[11][11],p[10][12]}), .w({r1[23][1],r1[22][4]})   ); 
    assign r1[22][5] = p[9][13];
    assign r1[22][6] = p[8][14];
    assign r1[22][7] = p[7][15]; //column 22
    
    FA e21(.p({p[15][8],p[14][9],p[13][10]}), .w({r1[24][0],r1[23][2]})   );
    assign r1[23][3] = p[12][11];
    assign r1[23][4] = p[11][12];
    assign r1[23][5] = p[10][13];
    assign r1[23][6] = p[9][14];
    assign r1[23][7] = p[8][15]; //column 23
    
    assign r1[24][1] = p[15][9];
    assign r1[24][2] = p[14][10];
    assign r1[24][3] = p[13][11];
    assign r1[24][4] = p[12][12];
    assign r1[24][5] = p[11][13];
    assign r1[24][6] = p[10][14];
    assign r1[24][7] = p[9][15]; //column 24
    
    assign r1[25][0] = p[15][10];
    assign r1[25][1] = p[14][11];
    assign r1[25][2] = p[13][12];
    assign r1[25][3] = p[12][13];
    assign r1[25][4] = p[11][14];
    assign r1[25][5] = p[10][15]; //column 25
    
    assign r1[26][0] = p[15][11];
    assign r1[26][1] = p[14][12];
    assign r1[26][2] = p[13][13];
    assign r1[26][3] = p[12][14];
    assign r1[26][4] = p[11][15]; //column 26
    
    assign r1[27][0] = p[15][12];
    assign r1[27][1] = p[14][13];
    assign r1[27][2] = p[13][14];
    assign r1[27][3] = p[12][15]; //column 27
    
    assign r1[28][0] = p[15][13];
    assign r1[28][1] = p[14][14];
    assign r1[28][2] = p[13][15]; //column 28
    
    assign r1[29][0] = p[15][14];
    assign r1[29][1] = p[14][15]; //column 29
   
    assign r1[30][0] = p[15][15]; //column 30
    
    ////////////////////////////////////////// PP REDUCTION STEP TWO   ////////////////////////  
    wire r2[30:0][3:0] ; // outputs of first reduction
    
    assign r2[0][0] = r1[0][0];// column 0
    
    assign r2[1][0] = r1[1][0];
    assign r2[1][1] = r1[1][1];// column 1
    
    assign r2[2][0] = r1[2][0];
    assign r2[2][1] = r1[2][1];// column 2
    
    assign r2[3][0] = r1[3][0];
    assign r2[3][1] = r1[3][1];// column 3
    
    compressor3_2 c16   (.p({r1[4][0]   ,r1[4][1]   ,r1[4][2]}),                                                       .w({r2[4][0]  ,r2[4][1]})); // column 4
    compressor3_2 c17   (.p({r1[5][0]   ,r1[5][1]   ,r1[5][2]}),                                                       .w({r2[5][0]  ,r2[5][1]})); // column 5
    compressor4_2 c18   (.p({r1[6][0]   ,r1[6][1]   ,r1[6][2]  ,r1[6][3]}),                                            .w({r2[6][0]  ,r2[6][1]})); // column 6
    compressor4_2 c19   (.p({r1[7][0]   ,r1[7][1]   ,r1[7][2]  ,r1[7][3]}),                                            .w({r2[7][0]  ,r2[7][1]})); // column 7
    compressor5_3 c20   (.p({r1[8][0]   ,r1[8][1]   ,r1[8][2]  ,r1[8][3]  ,r1[8][4]}),                                 .w({r2[8][0]  ,r2[8][1] ,r2[8][2]})); // column 8
    compressor5_3 c21   (.p({r1[9][0]   ,r1[9][1]   ,r1[9][2]  ,r1[9][3]  ,r1[9][4]}),                                 .w({r2[9][0]  ,r2[9][1] ,r2[9][2]})); // column 9
    compressor6_3 c22   (.p({r1[10][0]  ,r1[10][1]  ,r1[10][2] ,r1[10][3] ,r1[10][4],r1[10][5]}),                      .w({r2[10][0] ,r2[10][1],r2[10][2]})); // column 10
    compressor6_3 c23   (.p({r1[11][0]  ,r1[11][1]  ,r1[11][2] ,r1[11][3] ,r1[11][4],r1[11][5]}),                      .w({r2[11][0] ,r2[11][1],r2[11][2]})); // column 11
    compressor7_4 c24   (.p({r1[12][0]  ,r1[12][1]  ,r1[12][2] ,r1[12][3] ,r1[12][4],r1[12][5],r1[12][6]}),            .w({r2[12][0] ,r2[12][1],r2[12][2],r2[12][3]})); // column 12
    compressor7_4 c25   (.p({r1[13][0]  ,r1[13][1]  ,r1[13][2] ,r1[13][3] ,r1[13][4],r1[13][5],r1[13][6]}),            .w({r2[13][0] ,r2[13][1],r2[13][2],r2[13][3]})); // column 13
    compressor8_4 c26   (.p({r1[14][0]  ,r1[14][1]  ,r1[14][2] ,r1[14][3] ,r1[14][4],r1[14][5],r1[14][6],r1[14][7]}),  .w({r2[14][0] ,r2[14][1],r2[14][2],r2[14][3]})); // column 14
    compressor8_4 c27   (.p({r1[15][0]  ,r1[15][1]  ,r1[15][2] ,r1[15][3] ,r1[15][4],r1[15][5],r1[15][6],r1[15][7]}),  .w({r2[15][0] ,r2[15][1],r2[15][2],r2[15][3]})); // column 15
    compressor8_4 c28   (.p({r1[16][0]  ,r1[16][1]  ,r1[16][2] ,r1[16][3] ,r1[16][4],r1[16][5],r1[16][6],r1[16][7]}),  .w({r2[16][0] ,r2[16][1],r2[16][2],r2[16][3]})); // column 16
    compressor8_4 c29   (.p({r1[17][0]  ,r1[17][1]  ,r1[17][2] ,r1[17][3] ,r1[17][4],r1[17][5],r1[17][6],r1[17][7]}),  .w({r2[17][0] ,r2[17][1],r2[17][2],r2[17][3]})); // column 17
    compressor8_4 c30   (.p({r1[18][0]  ,r1[18][1]  ,r1[18][2] ,r1[18][3] ,r1[18][4],r1[18][5],r1[18][6],r1[18][7]}),  .w({r2[18][0] ,r2[18][1],r2[18][2],r2[18][3]})); // column 18
    compressor8_4 c31   (.p({r1[19][0]  ,r1[19][1]  ,r1[19][2] ,r1[19][3] ,r1[19][4],r1[19][5],r1[19][6],r1[19][7]}),  .w({r2[19][0] ,r2[19][1],r2[19][2],r2[19][3]})); // column 19
    compressor8_4 c32   (.p({r1[20][0]  ,r1[20][1]  ,r1[20][2] ,r1[20][3] ,r1[20][4],r1[20][5],r1[20][6],r1[20][7]}),  .w({r2[20][0] ,r2[20][1],r2[20][2],r2[20][3]})); // column 20
    compressor8_4 c33   (.p({r1[21][0]  ,r1[21][1]  ,r1[21][2] ,r1[21][3] ,r1[21][4],r1[21][5],r1[21][6],r1[21][7]}),  .w({r2[21][0] ,r2[21][1],r2[21][2],r2[21][3]})); // column 21
    compressor8_4 c34   (.p({r1[22][0]  ,r1[22][1]  ,r1[22][2] ,r1[22][3] ,r1[22][4],r1[22][5],r1[22][6],r1[22][7]}),  .w({r2[22][0] ,r2[22][1],r2[22][2],r2[22][3]})); // column 22
    compressor8_4 c35   (.p({r1[23][0]  ,r1[23][1]  ,r1[23][2] ,r1[23][3] ,r1[23][4],r1[23][5],r1[23][6],r1[23][7]}),  .w({r2[23][0] ,r2[23][1],r2[23][2],r2[23][3]})); // column 23
    
    FA e22(.p({r1[24][0],r1[24][1],r1[24][2]}), .w({r2[25][0],r2[24][0]})   );
    FA e23(.p({r1[24][3],r1[24][4],r1[24][5]}), .w({r2[25][1],r2[24][1]})   ); 
    assign r2[24][2] = r1[24][6];
    assign r2[24][3] = r1[24][7]; // column 24
    
    FA e24(.p({r1[25][0],r1[25][1],r1[25][2]}), .w({r2[26][0],r2[25][2]})   );
    FA e25(.p({r1[25][3],r1[25][4],r1[25][5]}), .w({r2[26][1],r2[25][3]})   ); // column 25
    
    FA e26(.p({r1[26][0],r1[26][1],r1[26][2]}), .w({r2[27][0],r2[26][2]})   );
    HA e27(.p({r1[26][3],r1[26][4]}),           .w({r2[27][1],r2[26][3]})   ); // column 26
    
    FA e28(.p({r1[27][0],r1[27][1],r1[27][2]}), .w({r2[28][0],r2[27][2]})   ); 
    assign r2[27][3] = r1[27][3]; // column 27
						
    assign r2[28][1] = r1[28][0];
    assign r2[28][2] = r1[28][1];
    assign r2[28][3] = r1[28][2]; //column 28
						
    assign r2[29][0] = r1[29][0];
    assign r2[29][1] = r1[29][1]; //column 29
						
    assign r2[30][0] = r1[30][0]; //column 30
    
    ////////////////////////////////////////// PP REDUCTION STEP THREE   ////////////////////////
	wire r3[30:0][1:0] ; // outputs of second reduction
	
	assign r3[0][0] = r2[0][0];// column 0
    
    assign r3[1][0] = r2[1][0];
    assign r3[1][1] = r2[1][1];// column 1
    
    assign r3[2][0] = r2[2][0];
    assign r3[2][1] = r2[2][1];// column 2
    
    assign r3[3][0] = r2[3][0];
    assign r3[3][1] = r2[3][1];// column 3
    
    assign r3[4][0] = r2[4][0];
    assign r3[4][1] = r2[4][1];// column 4
    
    assign r3[5][0] = r2[5][0];
    assign r3[5][1] = r2[5][1];// column 5
    
    assign r3[6][0] = r2[6][0];
    assign r3[6][1] = r2[6][1];// column 6
	
	assign r3[7][0] = r2[7][0];
    assign r3[7][1] = r2[7][1];// column 7

    compressor3_2 c36   (.p({r2[8][0]   ,r2[8][1]   ,r2[8][2]}),              .w({r3[8][0]   ,r3[8][1]})); // column 8
	compressor3_2 c37   (.p({r2[9][0]   ,r2[9][1]   ,r2[9][2]}),              .w({r3[9][0]   ,r3[9][1]})); // column 9
	compressor3_2 c38   (.p({r2[10][0]  ,r2[10][1]  ,r2[10][2]}),             .w({r3[10][0]  ,r3[10][1]})); // column 10
	compressor3_2 c39   (.p({r2[11][0]  ,r2[11][1]  ,r2[11][2]}),             .w({r3[11][0]  ,r3[11][1]})); // column 11
	compressor4_2 c40   (.p({r2[12][0]  ,r2[12][1]  ,r2[12][2] ,r2[12][3]}),  .w({r3[12][0]  ,r3[12][1]})); // column 12
	compressor4_2 c41   (.p({r2[13][0]  ,r2[13][1]  ,r2[13][2] ,r2[13][3]}),  .w({r3[13][0]  ,r3[13][1]})); // column 13
	compressor4_2 c42   (.p({r2[14][0]  ,r2[14][1]  ,r2[14][2] ,r2[14][3]}),  .w({r3[14][0]  ,r3[14][1]})); // column 14
	compressor4_2 c43   (.p({r2[15][0]  ,r2[15][1]  ,r2[15][2] ,r2[15][3]}),  .w({r3[15][0]  ,r3[15][1]})); // column 15
	compressor4_2 c44   (.p({r2[16][0]  ,r2[16][1]  ,r2[16][2] ,r2[16][3]}),  .w({r3[16][0]  ,r3[16][1]})); // column 16
	compressor4_2 c45   (.p({r2[17][0]  ,r2[17][1]  ,r2[17][2] ,r2[17][3]}),  .w({r3[17][0]  ,r3[17][1]})); // column 17
	compressor4_2 c46   (.p({r2[18][0]  ,r2[18][1]  ,r2[18][2] ,r2[18][3]}),  .w({r3[18][0]  ,r3[18][1]})); // column 18
	compressor4_2 c47   (.p({r2[19][0]  ,r2[19][1]  ,r2[19][2] ,r2[19][3]}),  .w({r3[19][0]  ,r3[19][1]})); // column 19
	compressor4_2 c48   (.p({r2[20][0]  ,r2[20][1]  ,r2[20][2] ,r2[20][3]}),  .w({r3[20][0]  ,r3[20][1]})); // column 20
	compressor4_2 c49   (.p({r2[21][0]  ,r2[21][1]  ,r2[21][2] ,r2[21][3]}),  .w({r3[21][0]  ,r3[21][1]})); // column 21
	compressor4_2 c51   (.p({r2[22][0]  ,r2[22][1]  ,r2[22][2] ,r2[22][3]}),  .w({r3[22][0]  ,r3[22][1]})); // column 22
	compressor4_2 c52   (.p({r2[23][0]  ,r2[23][1]  ,r2[23][2] ,r2[23][3]}),  .w({r3[23][0]  ,r3[23][1]})); // column 23
	compressor4_2 c53   (.p({r2[24][0]  ,r2[24][1]  ,r2[24][2] ,r2[24][3]}),  .w({r3[24][0]  ,r3[24][1]})); // column 24
	compressor4_2 c54   (.p({r2[25][0]  ,r2[25][1]  ,r2[25][2] ,r2[25][3]}),  .w({r3[25][0]  ,r3[25][1]})); // column 25
	compressor4_2 c55   (.p({r2[26][0]  ,r2[26][1]  ,r2[26][2] ,r2[26][3]}),  .w({r3[26][0]  ,r3[26][1]})); // column 26
	compressor4_2 c56   (.p({r2[27][0]  ,r2[27][1]  ,r2[27][2] ,r2[27][3]}),  .w({r3[27][0]  ,r3[27][1]})); // column 27
	                
	FA e29(.p({r2[28][0],r2[28][1],r2[28][2]}), .w({r3[29][0],r3[28][0]})   ); 
    assign r3[28][1] = r2[28][3]; // column 28
	
	HA e30(.p({r2[29][0],r2[29][1]}), .w({r3[30][0],r3[29][1]})   ); // column 29
	
    assign r3[30][1] = r2[30][0];// column 30
	
	assign r3[0][1] = 1'b0; // the third reduced pp doesnt provide value
	
	////////////////////////////////////////// Outputs of processing block   ////////////////////////
	assign out1[0] = r3[0][0];    
    assign out1[1] = r3[1][0];
    assign out1[2] = r3[2][0];
    assign out1[3] = r3[3][0];
    assign out1[4] = r3[4][0];
    assign out1[5] = r3[5][0];
    assign out1[6] = r3[6][0];
    assign out1[7] = r3[7][0];
    assign out1[8] = r3[8][0];
    assign out1[9] = r3[9][0];
    assign out1[10] = r3[10][0];
    assign out1[11] = r3[11][0];
    assign out1[12] = r3[12][0];
    assign out1[13] = r3[13][0];
    assign out1[14] = r3[14][0];
	assign out1[15] = r3[15][0];
    assign out1[16] = r3[16][0];
    assign out1[17] = r3[17][0];
    assign out1[18] = r3[18][0];
    assign out1[19] = r3[19][0];
	assign out1[20] = r3[20][0];
	assign out1[21] = r3[21][0];
    assign out1[22] = r3[22][0];
    assign out1[23] = r3[23][0];
    assign out1[24] = r3[24][0];
    assign out1[25] = r3[25][0];
    assign out1[26] = r3[26][0];
    assign out1[27] = r3[27][0];
    assign out1[28] = r3[28][0];
    assign out1[29] = r3[29][0];
    assign out1[30] = r3[30][0];
    
    assign out2[0] = r3[0][1];    
    assign out2[1] = r3[1][1];
    assign out2[2] = r3[2][1];
    assign out2[3] = r3[3][1];
    assign out2[4] = r3[4][1];
    assign out2[5] = r3[5][1];
    assign out2[6] = r3[6][1];
    assign out2[7] = r3[7][1];
    assign out2[8] = r3[8][1];
    assign out2[9] = r3[9][1];
    assign out2[10] = r3[10][1];
    assign out2[11] = r3[11][1];
    assign out2[12] = r3[12][1];
    assign out2[13] = r3[13][1];
    assign out2[14] = r3[14][1];
	assign out2[15] = r3[15][1];
    assign out2[16] = r3[16][1];
    assign out2[17] = r3[17][1];
    assign out2[18] = r3[18][1];
    assign out2[19] = r3[19][1];
	assign out2[20] = r3[20][1];
	assign out2[21] = r3[21][1];
    assign out2[22] = r3[22][1];
    assign out2[23] = r3[23][1];
    assign out2[24] = r3[24][1];
    assign out2[25] = r3[25][1];
    assign out2[26] = r3[26][1];
    assign out2[27] = r3[27][1];
    assign out2[28] = r3[28][1];
    assign out2[29] = r3[29][1];
    assign out2[30] = r3[30][1];
	
 endmodule 